library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity HttpServer is
  port (
    clk : in std_logic;
    reset : in std_logic;
    buffer_address : in signed(32-1 downto 0);
    buffer_we : in std_logic;
    buffer_oe : in std_logic;
    buffer_din : in signed(8-1 downto 0);
    buffer_dout : out signed(8-1 downto 0);
    buffer_length : out signed(32-1 downto 0);
    arg0_in : in signed(8-1 downto 0);
    arg0_we : in std_logic;
    arg0_out : out signed(8-1 downto 0);
    arg1_in : in signed(8-1 downto 0);
    arg1_we : in std_logic;
    arg1_out : out signed(8-1 downto 0);
    action_len : in signed(32-1 downto 0);
    init_contents_busy : out std_logic;
    init_contents_req : in std_logic;
    ready_contents_return : out signed(32-1 downto 0);
    ready_contents_busy : out std_logic;
    ready_contents_req : in std_logic;
    action_return : out signed(32-1 downto 0);
    action_busy : out std_logic;
    action_req : in std_logic
  );
end HttpServer;

architecture RTL of HttpServer is

  component http_response_header
    port (
      clk : in std_logic;
      reset : in std_logic;
      data_length : out signed(32-1 downto 0);
      data_address : in signed(32-1 downto 0);
      data_din : in signed(32-1 downto 0);
      data_dout : out signed(32-1 downto 0);
      data_we : in std_logic;
      data_oe : in std_logic;
      length : out signed(32-1 downto 0)
    );
  end component http_response_header;
  component dualportram
    generic (
      WIDTH : integer := 8;
      DEPTH : integer := 10;
      WORDS : integer := 1024
    );
    port (
      clk : in std_logic;
      reset : in std_logic;
      length : out signed(31 downto 0);
      address : in signed(31 downto 0);
      din : in signed(WIDTH-1 downto 0);
      dout : out signed(WIDTH-1 downto 0);
      we : in std_logic;
      oe : in std_logic;
      address_b : in signed(31 downto 0);
      din_b : in signed(WIDTH-1 downto 0);
      dout_b : out signed(WIDTH-1 downto 0);
      we_b : in std_logic;
      oe_b : in std_logic
    );
  end component dualportram;
  component singleportram
    generic (
      WIDTH : integer := 32;
      DEPTH : integer := 10;
      WORDS : integer := 1024
    );
    port (
      clk : in std_logic;
      reset : in std_logic;
      length : out signed(31 downto 0);
      address_b : in signed(31 downto 0);
      din_b : in signed(WIDTH-1 downto 0);
      dout_b : out signed(WIDTH-1 downto 0);
      we_b : in std_logic;
      oe_b : in std_logic
    );
  end component singleportram;
  component Misc
    port (
      clk : in std_logic;
      reset : in std_logic;
      quant_in : in signed(32-1 downto 0);
      quant_we : in std_logic;
      quant_out : out signed(32-1 downto 0);
      remainder_in : in signed(32-1 downto 0);
      remainder_we : in std_logic;
      remainder_out : out signed(32-1 downto 0);
      simple_div_n : in signed(32-1 downto 0);
      simple_div_d : in signed(32-1 downto 0);
      i_to_4digit_ascii_x : in signed(32-1 downto 0);
      i_to_4digit_ascii_flag : in std_logic;
      isHex_v : in signed(8-1 downto 0);
      toHex1_v : in signed(8-1 downto 0);
      toHex2_v0 : in signed(8-1 downto 0);
      toHex2_v1 : in signed(8-1 downto 0);
      simple_div_return : out signed(32-1 downto 0);
      simple_div_busy : out std_logic;
      simple_div_req : in std_logic;
      i_to_4digit_ascii_return : out signed(32-1 downto 0);
      i_to_4digit_ascii_busy : out std_logic;
      i_to_4digit_ascii_req : in std_logic;
      isHex_return : out std_logic;
      isHex_busy : out std_logic;
      isHex_req : in std_logic;
      toHex1_return : out signed(32-1 downto 0);
      toHex1_busy : out std_logic;
      toHex1_req : in std_logic;
      toHex2_return : out signed(32-1 downto 0);
      toHex2_busy : out std_logic;
      toHex2_req : in std_logic
    );
  end component Misc;

  signal clk_sig : std_logic;
  signal reset_sig : std_logic;
  signal buffer_address_sig : signed(32-1 downto 0);
  signal buffer_we_sig : std_logic;
  signal buffer_oe_sig : std_logic;
  signal buffer_din_sig : signed(8-1 downto 0);
  signal buffer_dout_sig : signed(8-1 downto 0);
  signal buffer_length_sig : signed(32-1 downto 0);
  signal arg0_in_sig : signed(8-1 downto 0);
  signal arg0_we_sig : std_logic;
  signal arg0_out_sig : signed(8-1 downto 0);
  signal arg1_in_sig : signed(8-1 downto 0);
  signal arg1_we_sig : std_logic;
  signal arg1_out_sig : signed(8-1 downto 0);
  signal action_len_sig : signed(32-1 downto 0);
  signal init_contents_busy_sig : std_logic := '1';
  signal init_contents_req_sig : std_logic;
  signal ready_contents_return_sig : signed(32-1 downto 0) := (others => '0');
  signal ready_contents_busy_sig : std_logic := '1';
  signal ready_contents_req_sig : std_logic;
  signal action_return_sig : signed(32-1 downto 0) := (others => '0');
  signal action_busy_sig : std_logic := '1';
  signal action_req_sig : std_logic;

  signal class_resp_0000_clk : std_logic;
  signal class_resp_0000_reset : std_logic;
  signal class_resp_0000_data_length : signed(32-1 downto 0);
  signal class_resp_0000_data_address : signed(32-1 downto 0) := (others => '0');
  signal class_resp_0000_data_din : signed(32-1 downto 0) := (others => '0');
  signal class_resp_0000_data_dout : signed(32-1 downto 0);
  signal class_resp_0000_data_we : std_logic := '0';
  signal class_resp_0000_data_oe : std_logic := '0';
  signal class_resp_0000_length : signed(32-1 downto 0);
  signal class_buffer_0002_clk : std_logic;
  signal class_buffer_0002_reset : std_logic;
  signal class_buffer_0002_length : signed(32-1 downto 0);
  signal class_buffer_0002_address : signed(32-1 downto 0);
  signal class_buffer_0002_din : signed(8-1 downto 0);
  signal class_buffer_0002_dout : signed(8-1 downto 0);
  signal class_buffer_0002_we : std_logic;
  signal class_buffer_0002_oe : std_logic;
  signal class_buffer_0002_address_b : signed(32-1 downto 0) := (others => '0');
  signal class_buffer_0002_din_b : signed(8-1 downto 0) := (others => '0');
  signal class_buffer_0002_dout_b : signed(8-1 downto 0);
  signal class_buffer_0002_we_b : std_logic := '0';
  signal class_buffer_0002_oe_b : std_logic := '0';
  signal class_data_0003_clk : std_logic;
  signal class_data_0003_reset : std_logic;
  signal class_data_0003_length : signed(32-1 downto 0);
  signal class_data_0003_address_b : signed(32-1 downto 0) := (others => '0');
  signal class_data_0003_din_b : signed(32-1 downto 0) := (others => '0');
  signal class_data_0003_dout_b : signed(32-1 downto 0);
  signal class_data_0003_we_b : std_logic := '0';
  signal class_data_0003_oe_b : std_logic := '0';
  signal class_content_words_0004 : signed(32-1 downto 0) := X"00000008";
  signal class_content_length_field_0_0005 : signed(32-1 downto 0) := (others => '0');
  signal class_content_length_field_1_0006 : signed(32-1 downto 0) := (others => '0');
  signal class_content_length_field_2_0007 : signed(32-1 downto 0) := (others => '0');
  signal class_misc_0008_clk : std_logic;
  signal class_misc_0008_reset : std_logic;
  signal class_misc_0008_quant_in : signed(32-1 downto 0) := (others => '0');
  signal class_misc_0008_quant_we : std_logic := '0';
  signal class_misc_0008_quant_out : signed(32-1 downto 0);
  signal class_misc_0008_remainder_in : signed(32-1 downto 0) := (others => '0');
  signal class_misc_0008_remainder_we : std_logic := '0';
  signal class_misc_0008_remainder_out : signed(32-1 downto 0);
  signal class_misc_0008_simple_div_n : signed(32-1 downto 0) := (others => '0');
  signal class_misc_0008_simple_div_d : signed(32-1 downto 0) := (others => '0');
  signal class_misc_0008_i_to_4digit_ascii_x : signed(32-1 downto 0) := (others => '0');
  signal class_misc_0008_i_to_4digit_ascii_flag : std_logic := '0';
  signal class_misc_0008_isHex_v : signed(8-1 downto 0) := (others => '0');
  signal class_misc_0008_toHex1_v : signed(8-1 downto 0) := (others => '0');
  signal class_misc_0008_toHex2_v0 : signed(8-1 downto 0) := (others => '0');
  signal class_misc_0008_toHex2_v1 : signed(8-1 downto 0) := (others => '0');
  signal class_misc_0008_simple_div_return : signed(32-1 downto 0);
  signal class_misc_0008_simple_div_busy : std_logic;
  signal class_misc_0008_simple_div_req : std_logic := '0';
  signal class_misc_0008_i_to_4digit_ascii_return : signed(32-1 downto 0);
  signal class_misc_0008_i_to_4digit_ascii_busy : std_logic;
  signal class_misc_0008_i_to_4digit_ascii_req : std_logic := '0';
  signal class_misc_0008_isHex_return : std_logic;
  signal class_misc_0008_isHex_busy : std_logic;
  signal class_misc_0008_isHex_req : std_logic := '0';
  signal class_misc_0008_toHex1_return : signed(32-1 downto 0);
  signal class_misc_0008_toHex1_busy : std_logic;
  signal class_misc_0008_toHex1_req : std_logic := '0';
  signal class_misc_0008_toHex2_return : signed(32-1 downto 0);
  signal class_misc_0008_toHex2_busy : std_logic;
  signal class_misc_0008_toHex2_req : std_logic := '0';
  signal class_arg0_0010 : signed(8-1 downto 0) := X"20";
  signal class_arg0_0010_mux : signed(8-1 downto 0);
  signal tmp_0001 : signed(8-1 downto 0);
  signal class_arg1_0011 : signed(8-1 downto 0) := X"20";
  signal class_arg1_0011_mux : signed(8-1 downto 0);
  signal tmp_0002 : signed(8-1 downto 0);
  signal pack_a_0012 : std_logic_vector(16-1 downto 0) := (others => '0');
  signal pack_a_local : std_logic_vector(16-1 downto 0) := (others => '0');
  signal pack_b_0013 : std_logic_vector(16-1 downto 0) := (others => '0');
  signal pack_b_local : std_logic_vector(16-1 downto 0) := (others => '0');
  signal pack_c_0014 : std_logic_vector(16-1 downto 0) := (others => '0');
  signal pack_c_local : std_logic_vector(16-1 downto 0) := (others => '0');
  signal pack_d_0015 : std_logic_vector(16-1 downto 0) := (others => '0');
  signal pack_d_local : std_logic_vector(16-1 downto 0) := (others => '0');
  signal cast_expr_00016 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00017 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00018 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00019 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00020 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00021 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00022 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00023 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00024 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00025 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00026 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00027 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00028 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00029 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00030 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00031 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00032 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00033 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00034 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00035 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00036 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00037 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00038 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00039 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00040 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00041 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00042 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00043 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00044 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00045 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00046 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00047 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00048 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00049 : signed(32-1 downto 0) := (others => '0');
  signal init_contents_v_0050 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00051 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00052 : signed(32-1 downto 0) := (others => '0');
  signal init_contents_bytes_2_0053 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00054 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00055 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00056 : signed(32-1 downto 0) := (others => '0');
  signal init_contents_bytes_1_0057 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00058 : signed(32-1 downto 0) := (others => '0');
  signal init_contents_bytes_0_0059 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00060 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00061 : std_logic := '0';
  signal method_result_00062 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00063 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00064 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00065 : std_logic := '0';
  signal method_result_00066 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00067 : signed(32-1 downto 0) := (others => '0');
  signal method_result_00068 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00096 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00097 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00098 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00099 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00100 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00101 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00102 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00103 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00104 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00105 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00106 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00107 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00108 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00109 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00110 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00111 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00112 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00113 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00114 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00115 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00116 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00117 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00118 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00119 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00120 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00121 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00122 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00123 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00124 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00125 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00126 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00127 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00128 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00129 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00130 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00131 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00132 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00133 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00134 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00135 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00136 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00137 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00138 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00139 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00140 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00141 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00142 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00143 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00144 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00145 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00146 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00147 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00148 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00149 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00150 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00151 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00152 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00153 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00154 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00155 : signed(8-1 downto 0) := (others => '0');
  signal ready_contents_offset_0156 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00157 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00187 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00188 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00189 : signed(32-1 downto 0) := (others => '0');
  signal ready_contents_i_0069 : signed(32-1 downto 0) := X"00000000";
  signal field_access_00070 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00071 : std_logic := '0';
  signal unary_expr_00072 : signed(32-1 downto 0) := (others => '0');
  signal ready_contents_v_0073 : signed(32-1 downto 0) := (others => '0');
  signal field_access_00074 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00075 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00076 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00077 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00078 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00079 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00080 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00081 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00082 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00083 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00084 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00085 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00086 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00087 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00088 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00089 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00090 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00091 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00092 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00093 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00094 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00095 : signed(8-1 downto 0) := (others => '0');
  signal ready_contents_i_0158 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00159 : std_logic := '0';
  signal unary_expr_00160 : signed(32-1 downto 0) := (others => '0');
  signal ready_contents_v_0161 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00162 : signed(32-1 downto 0) := (others => '0');
  signal ready_contents_ptr_0163 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00164 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00165 : signed(32-1 downto 0) := (others => '0');
  signal binary_expr_00166 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00167 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00168 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00169 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00170 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00171 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00172 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00173 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00174 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00175 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00176 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00177 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00178 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00179 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00180 : signed(32-1 downto 0) := (others => '0');
  signal cast_expr_00181 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00182 : std_logic := '0';
  signal binary_expr_00183 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00184 : signed(8-1 downto 0) := (others => '0');
  signal binary_expr_00185 : signed(32-1 downto 0) := (others => '0');
  signal array_access_00186 : signed(8-1 downto 0) := (others => '0');
  signal action_len_0190 : signed(32-1 downto 0) := (others => '0');
  signal action_len_local : signed(32-1 downto 0) := (others => '0');
  signal action_S_0191 : signed(32-1 downto 0) := X"00000000";
  signal action_v0_0192 : signed(8-1 downto 0) := X"00";
  signal action_v1_0193 : signed(8-1 downto 0) := X"00";
  signal action_v_0204 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00205 : std_logic := '0';
  signal action_i_0194 : signed(32-1 downto 0) := X"00000000";
  signal binary_expr_00195 : std_logic := '0';
  signal unary_expr_00196 : signed(32-1 downto 0) := (others => '0');
  signal action_b_0197 : signed(8-1 downto 0) := (others => '0');
  signal array_access_00198 : signed(8-1 downto 0) := (others => '0');
  signal method_result_00199 : std_logic := '0';
  signal method_result_00200 : std_logic := '0';
  signal binary_expr_00201 : std_logic := '0';
  signal binary_expr_00202 : std_logic := '0';
  signal binary_expr_00203 : std_logic := '0';
  signal method_result_00206 : signed(32-1 downto 0) := (others => '0');
  signal pack_return : signed(32-1 downto 0) := (others => '0');
  signal pack_busy : std_logic := '0';
  signal pack_req_flag : std_logic;
  signal pack_req_local : std_logic := '0';
  signal init_contents_req_flag : std_logic;
  signal init_contents_req_local : std_logic := '0';
  signal tmp_0003 : std_logic;
  signal ready_contents_req_flag : std_logic;
  signal ready_contents_req_local : std_logic := '0';
  signal tmp_0004 : std_logic;
  signal action_req_flag : std_logic;
  signal action_req_local : std_logic := '0';
  signal tmp_0005 : std_logic;
  type Type_pack_method is (
    pack_method_IDLE,
    pack_method_S_0000,
    pack_method_S_0001,
    pack_method_S_0002,
    pack_method_S_0016,
    pack_method_S_0017  
  );
  signal pack_method : Type_pack_method := pack_method_IDLE;
  signal pack_method_delay : signed(32-1 downto 0) := (others => '0');
  signal pack_req_flag_d : std_logic := '0';
  signal pack_req_flag_edge : std_logic;
  signal tmp_0006 : std_logic;
  signal tmp_0007 : std_logic;
  signal tmp_0008 : std_logic;
  signal tmp_0009 : std_logic;
  signal tmp_0010 : std_logic;
  signal tmp_0011 : std_logic;
  signal tmp_0012 : std_logic;
  signal tmp_0013 : std_logic;
  signal tmp_0014 : std_logic_vector(32-1 downto 0);
  signal tmp_0015 : std_logic_vector(32-1 downto 0);
  signal tmp_0016 : std_logic_vector(32-1 downto 0);
  signal tmp_0017 : std_logic_vector(32-1 downto 0);
  signal tmp_0018 : signed(32-1 downto 0);
  signal tmp_0019 : signed(32-1 downto 0);
  signal tmp_0020 : signed(32-1 downto 0);
  signal tmp_0021 : signed(32-1 downto 0);
  signal tmp_0022 : signed(32-1 downto 0);
  signal tmp_0023 : signed(32-1 downto 0);
  signal tmp_0024 : signed(32-1 downto 0);
  signal tmp_0025 : signed(32-1 downto 0);
  signal tmp_0026 : signed(32-1 downto 0);
  signal tmp_0027 : signed(32-1 downto 0);
  type Type_init_contents_method is (
    init_contents_method_IDLE,
    init_contents_method_S_0000,
    init_contents_method_S_0001,
    init_contents_method_S_0002,
    init_contents_method_S_0003,
    init_contents_method_S_0004,
    init_contents_method_S_0005,
    init_contents_method_S_0006,
    init_contents_method_S_0007,
    init_contents_method_S_0008,
    init_contents_method_S_0009,
    init_contents_method_S_0010,
    init_contents_method_S_0011,
    init_contents_method_S_0012,
    init_contents_method_S_0013,
    init_contents_method_S_0014,
    init_contents_method_S_0015,
    init_contents_method_S_0016,
    init_contents_method_S_0017,
    init_contents_method_S_0018,
    init_contents_method_S_0019,
    init_contents_method_S_0020,
    init_contents_method_S_0021,
    init_contents_method_S_0022,
    init_contents_method_S_0023,
    init_contents_method_S_0024,
    init_contents_method_S_0025,
    init_contents_method_S_0026,
    init_contents_method_S_0027,
    init_contents_method_S_0028,
    init_contents_method_S_0029,
    init_contents_method_S_0030,
    init_contents_method_S_0031,
    init_contents_method_S_0035,
    init_contents_method_S_0036,
    init_contents_method_S_0037,
    init_contents_method_S_0038,
    init_contents_method_S_0039,
    init_contents_method_S_0040,
    init_contents_method_S_0041,
    init_contents_method_S_0042,
    init_contents_method_S_0043,
    init_contents_method_S_0044,
    init_contents_method_S_0046,
    init_contents_method_S_0047,
    init_contents_method_S_0048,
    init_contents_method_S_0049,
    init_contents_method_S_0050,
    init_contents_method_S_0051,
    init_contents_method_S_0052,
    init_contents_method_S_0053,
    init_contents_method_S_0054,
    init_contents_method_S_0055,
    init_contents_method_S_0056,
    init_contents_method_S_0057,
    init_contents_method_S_0058,
    init_contents_method_S_0059,
    init_contents_method_S_0060,
    init_contents_method_S_0061,
    init_contents_method_S_0062,
    init_contents_method_S_0063,
    init_contents_method_S_0064,
    init_contents_method_S_0066,
    init_contents_method_S_0067,
    init_contents_method_S_0068,
    init_contents_method_S_0069,
    init_contents_method_S_0070,
    init_contents_method_S_0003_body,
    init_contents_method_S_0003_wait,
    init_contents_method_S_0006_body,
    init_contents_method_S_0006_wait,
    init_contents_method_S_0009_body,
    init_contents_method_S_0009_wait,
    init_contents_method_S_0012_body,
    init_contents_method_S_0012_wait,
    init_contents_method_S_0015_body,
    init_contents_method_S_0015_wait,
    init_contents_method_S_0018_body,
    init_contents_method_S_0018_wait,
    init_contents_method_S_0021_body,
    init_contents_method_S_0021_wait,
    init_contents_method_S_0024_body,
    init_contents_method_S_0024_wait,
    init_contents_method_S_0027_body,
    init_contents_method_S_0027_wait,
    init_contents_method_S_0030_body,
    init_contents_method_S_0030_wait,
    init_contents_method_S_0035_body,
    init_contents_method_S_0035_wait,
    init_contents_method_S_0040_body,
    init_contents_method_S_0040_wait,
    init_contents_method_S_0048_body,
    init_contents_method_S_0048_wait,
    init_contents_method_S_0050_body,
    init_contents_method_S_0050_wait,
    init_contents_method_S_0052_body,
    init_contents_method_S_0052_wait,
    init_contents_method_S_0059_body,
    init_contents_method_S_0059_wait,
    init_contents_method_S_0061_body,
    init_contents_method_S_0061_wait,
    init_contents_method_S_0066_body,
    init_contents_method_S_0066_wait  
  );
  signal init_contents_method : Type_init_contents_method := init_contents_method_IDLE;
  signal init_contents_method_delay : signed(32-1 downto 0) := (others => '0');
  signal init_contents_req_flag_d : std_logic := '0';
  signal init_contents_req_flag_edge : std_logic;
  signal tmp_0028 : std_logic;
  signal tmp_0029 : std_logic;
  signal tmp_0030 : std_logic;
  signal tmp_0031 : std_logic;
  signal pack_call_flag_0003 : std_logic;
  signal tmp_0032 : std_logic;
  signal tmp_0033 : std_logic;
  signal tmp_0034 : std_logic;
  signal tmp_0035 : std_logic;
  signal pack_call_flag_0006 : std_logic;
  signal tmp_0036 : std_logic;
  signal tmp_0037 : std_logic;
  signal tmp_0038 : std_logic;
  signal tmp_0039 : std_logic;
  signal pack_call_flag_0009 : std_logic;
  signal tmp_0040 : std_logic;
  signal tmp_0041 : std_logic;
  signal tmp_0042 : std_logic;
  signal tmp_0043 : std_logic;
  signal pack_call_flag_0012 : std_logic;
  signal tmp_0044 : std_logic;
  signal tmp_0045 : std_logic;
  signal tmp_0046 : std_logic;
  signal tmp_0047 : std_logic;
  signal pack_call_flag_0015 : std_logic;
  signal tmp_0048 : std_logic;
  signal tmp_0049 : std_logic;
  signal tmp_0050 : std_logic;
  signal tmp_0051 : std_logic;
  signal pack_call_flag_0018 : std_logic;
  signal tmp_0052 : std_logic;
  signal tmp_0053 : std_logic;
  signal tmp_0054 : std_logic;
  signal tmp_0055 : std_logic;
  signal pack_call_flag_0021 : std_logic;
  signal tmp_0056 : std_logic;
  signal tmp_0057 : std_logic;
  signal tmp_0058 : std_logic;
  signal tmp_0059 : std_logic;
  signal pack_call_flag_0024 : std_logic;
  signal tmp_0060 : std_logic;
  signal tmp_0061 : std_logic;
  signal tmp_0062 : std_logic;
  signal tmp_0063 : std_logic;
  signal pack_call_flag_0027 : std_logic;
  signal tmp_0064 : std_logic;
  signal tmp_0065 : std_logic;
  signal tmp_0066 : std_logic;
  signal tmp_0067 : std_logic;
  signal pack_call_flag_0030 : std_logic;
  signal tmp_0068 : std_logic;
  signal tmp_0069 : std_logic;
  signal tmp_0070 : std_logic;
  signal tmp_0071 : std_logic;
  signal simple_div_ext_call_flag_0035 : std_logic;
  signal tmp_0072 : std_logic;
  signal tmp_0073 : std_logic;
  signal tmp_0074 : std_logic;
  signal tmp_0075 : std_logic;
  signal simple_div_ext_call_flag_0040 : std_logic;
  signal tmp_0076 : std_logic;
  signal tmp_0077 : std_logic;
  signal tmp_0078 : std_logic;
  signal tmp_0079 : std_logic;
  signal tmp_0080 : std_logic;
  signal tmp_0081 : std_logic;
  signal i_to_4digit_ascii_ext_call_flag_0048 : std_logic;
  signal tmp_0082 : std_logic;
  signal tmp_0083 : std_logic;
  signal tmp_0084 : std_logic;
  signal tmp_0085 : std_logic;
  signal i_to_4digit_ascii_ext_call_flag_0050 : std_logic;
  signal tmp_0086 : std_logic;
  signal tmp_0087 : std_logic;
  signal tmp_0088 : std_logic;
  signal tmp_0089 : std_logic;
  signal i_to_4digit_ascii_ext_call_flag_0052 : std_logic;
  signal tmp_0090 : std_logic;
  signal tmp_0091 : std_logic;
  signal tmp_0092 : std_logic;
  signal tmp_0093 : std_logic;
  signal tmp_0094 : std_logic;
  signal tmp_0095 : std_logic;
  signal i_to_4digit_ascii_ext_call_flag_0059 : std_logic;
  signal tmp_0096 : std_logic;
  signal tmp_0097 : std_logic;
  signal tmp_0098 : std_logic;
  signal tmp_0099 : std_logic;
  signal i_to_4digit_ascii_ext_call_flag_0061 : std_logic;
  signal tmp_0100 : std_logic;
  signal tmp_0101 : std_logic;
  signal tmp_0102 : std_logic;
  signal tmp_0103 : std_logic;
  signal i_to_4digit_ascii_ext_call_flag_0066 : std_logic;
  signal tmp_0104 : std_logic;
  signal tmp_0105 : std_logic;
  signal tmp_0106 : std_logic;
  signal tmp_0107 : std_logic;
  signal tmp_0108 : std_logic;
  signal tmp_0109 : std_logic;
  signal tmp_0110 : std_logic;
  signal tmp_0111 : std_logic;
  signal tmp_0112 : signed(32-1 downto 0);
  signal tmp_0113 : std_logic;
  signal tmp_0114 : std_logic;
  type Type_ready_contents_method is (
    ready_contents_method_IDLE,
    ready_contents_method_S_0000,
    ready_contents_method_S_0001,
    ready_contents_method_S_0002,
    ready_contents_method_S_0003,
    ready_contents_method_S_0004,
    ready_contents_method_S_0005,
    ready_contents_method_S_0006,
    ready_contents_method_S_0007,
    ready_contents_method_S_0009,
    ready_contents_method_S_0010,
    ready_contents_method_S_0011,
    ready_contents_method_S_0012,
    ready_contents_method_S_0015,
    ready_contents_method_S_0016,
    ready_contents_method_S_0021,
    ready_contents_method_S_0022,
    ready_contents_method_S_0027,
    ready_contents_method_S_0028,
    ready_contents_method_S_0033,
    ready_contents_method_S_0034,
    ready_contents_method_S_0037,
    ready_contents_method_S_0038,
    ready_contents_method_S_0040,
    ready_contents_method_S_0041,
    ready_contents_method_S_0046,
    ready_contents_method_S_0047,
    ready_contents_method_S_0052,
    ready_contents_method_S_0053,
    ready_contents_method_S_0058,
    ready_contents_method_S_0059,
    ready_contents_method_S_0064,
    ready_contents_method_S_0065,
    ready_contents_method_S_0070,
    ready_contents_method_S_0071,
    ready_contents_method_S_0076,
    ready_contents_method_S_0077,
    ready_contents_method_S_0082,
    ready_contents_method_S_0083,
    ready_contents_method_S_0088,
    ready_contents_method_S_0089,
    ready_contents_method_S_0094,
    ready_contents_method_S_0095,
    ready_contents_method_S_0100,
    ready_contents_method_S_0101,
    ready_contents_method_S_0106,
    ready_contents_method_S_0107,
    ready_contents_method_S_0110,
    ready_contents_method_S_0111,
    ready_contents_method_S_0113,
    ready_contents_method_S_0114,
    ready_contents_method_S_0115,
    ready_contents_method_S_0116,
    ready_contents_method_S_0118,
    ready_contents_method_S_0119,
    ready_contents_method_S_0120,
    ready_contents_method_S_0125,
    ready_contents_method_S_0126,
    ready_contents_method_S_0130,
    ready_contents_method_S_0131,
    ready_contents_method_S_0135,
    ready_contents_method_S_0136,
    ready_contents_method_S_0140,
    ready_contents_method_S_0141,
    ready_contents_method_S_0145,
    ready_contents_method_S_0146,
    ready_contents_method_S_0147,
    ready_contents_method_S_0148,
    ready_contents_method_S_0150,
    ready_contents_method_S_0151,
    ready_contents_method_S_0153,
    ready_contents_method_S_0154,
    ready_contents_method_S_0155,
    ready_contents_method_S_0156,
    ready_contents_method_S_0158,
    ready_contents_method_S_0159  
  );
  signal ready_contents_method : Type_ready_contents_method := ready_contents_method_IDLE;
  signal ready_contents_method_delay : signed(32-1 downto 0) := (others => '0');
  signal ready_contents_req_flag_d : std_logic := '0';
  signal ready_contents_req_flag_edge : std_logic;
  signal tmp_0115 : std_logic;
  signal tmp_0116 : std_logic;
  signal tmp_0117 : std_logic;
  signal tmp_0118 : std_logic;
  signal tmp_0119 : std_logic;
  signal tmp_0120 : std_logic;
  signal tmp_0121 : std_logic;
  signal tmp_0122 : std_logic;
  signal tmp_0123 : std_logic;
  signal tmp_0124 : std_logic;
  signal tmp_0125 : std_logic;
  signal tmp_0126 : std_logic;
  signal tmp_0127 : std_logic;
  signal tmp_0128 : std_logic;
  signal tmp_0129 : std_logic;
  signal tmp_0130 : signed(32-1 downto 0);
  signal tmp_0131 : signed(32-1 downto 0);
  signal tmp_0132 : signed(32-1 downto 0);
  signal tmp_0133 : signed(32-1 downto 0);
  signal tmp_0134 : signed(32-1 downto 0);
  signal tmp_0135 : signed(8-1 downto 0);
  signal tmp_0136 : signed(32-1 downto 0);
  signal tmp_0137 : signed(32-1 downto 0);
  signal tmp_0138 : signed(32-1 downto 0);
  signal tmp_0139 : signed(8-1 downto 0);
  signal tmp_0140 : signed(32-1 downto 0);
  signal tmp_0141 : signed(32-1 downto 0);
  signal tmp_0142 : signed(32-1 downto 0);
  signal tmp_0143 : signed(8-1 downto 0);
  signal tmp_0144 : signed(32-1 downto 0);
  signal tmp_0145 : signed(32-1 downto 0);
  signal tmp_0146 : signed(8-1 downto 0);
  signal tmp_0147 : signed(32-1 downto 0);
  signal tmp_0148 : signed(32-1 downto 0);
  signal tmp_0149 : signed(32-1 downto 0);
  signal tmp_0150 : signed(32-1 downto 0);
  signal tmp_0151 : signed(8-1 downto 0);
  signal tmp_0152 : signed(32-1 downto 0);
  signal tmp_0153 : signed(32-1 downto 0);
  signal tmp_0154 : signed(32-1 downto 0);
  signal tmp_0155 : signed(8-1 downto 0);
  signal tmp_0156 : signed(32-1 downto 0);
  signal tmp_0157 : signed(32-1 downto 0);
  signal tmp_0158 : signed(32-1 downto 0);
  signal tmp_0159 : signed(8-1 downto 0);
  signal tmp_0160 : signed(32-1 downto 0);
  signal tmp_0161 : signed(32-1 downto 0);
  signal tmp_0162 : signed(32-1 downto 0);
  signal tmp_0163 : signed(8-1 downto 0);
  signal tmp_0164 : signed(32-1 downto 0);
  signal tmp_0165 : signed(32-1 downto 0);
  signal tmp_0166 : signed(32-1 downto 0);
  signal tmp_0167 : signed(8-1 downto 0);
  signal tmp_0168 : signed(32-1 downto 0);
  signal tmp_0169 : signed(32-1 downto 0);
  signal tmp_0170 : signed(32-1 downto 0);
  signal tmp_0171 : signed(8-1 downto 0);
  signal tmp_0172 : signed(32-1 downto 0);
  signal tmp_0173 : signed(32-1 downto 0);
  signal tmp_0174 : signed(32-1 downto 0);
  signal tmp_0175 : signed(8-1 downto 0);
  signal tmp_0176 : signed(32-1 downto 0);
  signal tmp_0177 : signed(32-1 downto 0);
  signal tmp_0178 : signed(32-1 downto 0);
  signal tmp_0179 : signed(8-1 downto 0);
  signal tmp_0180 : signed(32-1 downto 0);
  signal tmp_0181 : signed(32-1 downto 0);
  signal tmp_0182 : signed(32-1 downto 0);
  signal tmp_0183 : signed(8-1 downto 0);
  signal tmp_0184 : signed(32-1 downto 0);
  signal tmp_0185 : signed(32-1 downto 0);
  signal tmp_0186 : signed(32-1 downto 0);
  signal tmp_0187 : signed(8-1 downto 0);
  signal tmp_0188 : signed(32-1 downto 0);
  signal tmp_0189 : signed(32-1 downto 0);
  signal tmp_0190 : signed(32-1 downto 0);
  signal tmp_0191 : signed(8-1 downto 0);
  signal tmp_0192 : signed(32-1 downto 0);
  signal tmp_0193 : signed(32-1 downto 0);
  signal tmp_0194 : signed(8-1 downto 0);
  signal tmp_0195 : std_logic;
  signal tmp_0196 : signed(32-1 downto 0);
  signal tmp_0197 : signed(32-1 downto 0);
  signal tmp_0198 : signed(32-1 downto 0);
  signal tmp_0199 : signed(32-1 downto 0);
  signal tmp_0200 : signed(32-1 downto 0);
  signal tmp_0201 : signed(32-1 downto 0);
  signal tmp_0202 : signed(8-1 downto 0);
  signal tmp_0203 : signed(32-1 downto 0);
  signal tmp_0204 : signed(32-1 downto 0);
  signal tmp_0205 : signed(8-1 downto 0);
  signal tmp_0206 : signed(32-1 downto 0);
  signal tmp_0207 : signed(32-1 downto 0);
  signal tmp_0208 : signed(8-1 downto 0);
  signal tmp_0209 : signed(32-1 downto 0);
  signal tmp_0210 : std_logic;
  signal tmp_0211 : signed(8-1 downto 0);
  signal tmp_0212 : signed(32-1 downto 0);
  signal tmp_0213 : signed(32-1 downto 0);
  signal tmp_0214 : signed(32-1 downto 0);
  signal tmp_0215 : signed(32-1 downto 0);
  type Type_action_method is (
    action_method_IDLE,
    action_method_S_0000,
    action_method_S_0001,
    action_method_S_0002,
    action_method_S_0006,
    action_method_S_0007,
    action_method_S_0008,
    action_method_S_0009,
    action_method_S_0011,
    action_method_S_0012,
    action_method_S_0013,
    action_method_S_0014,
    action_method_S_0015,
    action_method_S_0016,
    action_method_S_0017,
    action_method_S_0018,
    action_method_S_0019,
    action_method_S_0020,
    action_method_S_0021,
    action_method_S_0022,
    action_method_S_0023,
    action_method_S_0025,
    action_method_S_0026,
    action_method_S_0027,
    action_method_S_0028,
    action_method_S_0029,
    action_method_S_0030,
    action_method_S_0031,
    action_method_S_0032,
    action_method_S_0033,
    action_method_S_0035,
    action_method_S_0036,
    action_method_S_0037,
    action_method_S_0038,
    action_method_S_0039,
    action_method_S_0040,
    action_method_S_0041,
    action_method_S_0042,
    action_method_S_0043,
    action_method_S_0044,
    action_method_S_0045,
    action_method_S_0046,
    action_method_S_0047,
    action_method_S_0048,
    action_method_S_0049,
    action_method_S_0050,
    action_method_S_0051,
    action_method_S_0052,
    action_method_S_0053,
    action_method_S_0054,
    action_method_S_0055,
    action_method_S_0056,
    action_method_S_0057,
    action_method_S_0058,
    action_method_S_0059,
    action_method_S_0060,
    action_method_S_0061,
    action_method_S_0062,
    action_method_S_0063,
    action_method_S_0064,
    action_method_S_0065,
    action_method_S_0066,
    action_method_S_0067,
    action_method_S_0068,
    action_method_S_0070,
    action_method_S_0071,
    action_method_S_0072,
    action_method_S_0073,
    action_method_S_0076,
    action_method_S_0077,
    action_method_S_0079,
    action_method_S_0080,
    action_method_S_0081,
    action_method_S_0020_body,
    action_method_S_0020_wait,
    action_method_S_0030_body,
    action_method_S_0030_wait,
    action_method_S_0072_body,
    action_method_S_0072_wait  
  );
  signal action_method : Type_action_method := action_method_IDLE;
  signal action_method_delay : signed(32-1 downto 0) := (others => '0');
  signal action_req_flag_d : std_logic := '0';
  signal action_req_flag_edge : std_logic;
  signal tmp_0216 : std_logic;
  signal tmp_0217 : std_logic;
  signal tmp_0218 : std_logic;
  signal tmp_0219 : std_logic;
  signal tmp_0220 : std_logic;
  signal tmp_0221 : std_logic;
  signal tmp_0222 : std_logic;
  signal tmp_0223 : std_logic;
  signal tmp_0224 : std_logic;
  signal tmp_0225 : std_logic;
  signal tmp_0226 : std_logic;
  signal tmp_0227 : std_logic;
  signal isHex_ext_call_flag_0020 : std_logic;
  signal tmp_0228 : std_logic;
  signal tmp_0229 : std_logic;
  signal tmp_0230 : std_logic;
  signal tmp_0231 : std_logic;
  signal tmp_0232 : std_logic;
  signal tmp_0233 : std_logic;
  signal isHex_ext_call_flag_0030 : std_logic;
  signal tmp_0234 : std_logic;
  signal tmp_0235 : std_logic;
  signal tmp_0236 : std_logic;
  signal tmp_0237 : std_logic;
  signal tmp_0238 : std_logic;
  signal tmp_0239 : std_logic;
  signal tmp_0240 : std_logic;
  signal tmp_0241 : std_logic;
  signal tmp_0242 : std_logic;
  signal tmp_0243 : std_logic;
  signal tmp_0244 : std_logic;
  signal tmp_0245 : std_logic;
  signal tmp_0246 : std_logic;
  signal tmp_0247 : std_logic;
  signal toHex2_ext_call_flag_0072 : std_logic;
  signal tmp_0248 : std_logic;
  signal tmp_0249 : std_logic;
  signal tmp_0250 : std_logic;
  signal tmp_0251 : std_logic;
  signal tmp_0252 : std_logic;
  signal tmp_0253 : std_logic;
  signal tmp_0254 : std_logic;
  signal tmp_0255 : std_logic;
  signal tmp_0256 : signed(32-1 downto 0);
  signal tmp_0257 : std_logic;
  signal tmp_0258 : signed(32-1 downto 0);
  signal tmp_0259 : std_logic;
  signal tmp_0260 : std_logic;
  signal tmp_0261 : std_logic;
  signal tmp_0262 : std_logic;

begin

  clk_sig <= clk;
  reset_sig <= reset;
  buffer_address_sig <= buffer_address;
  buffer_we_sig <= buffer_we;
  buffer_oe_sig <= buffer_oe;
  buffer_din_sig <= buffer_din;
  buffer_dout <= buffer_dout_sig;
  buffer_dout_sig <= class_buffer_0002_dout;

  buffer_length <= buffer_length_sig;
  buffer_length_sig <= class_buffer_0002_length;

  arg0_in_sig <= arg0_in;
  arg0_we_sig <= arg0_we;
  arg0_out <= arg0_out_sig;
  arg0_out_sig <= class_arg0_0010;

  arg1_in_sig <= arg1_in;
  arg1_we_sig <= arg1_we;
  arg1_out <= arg1_out_sig;
  arg1_out_sig <= class_arg1_0011;

  action_len_sig <= action_len;
  init_contents_busy <= init_contents_busy_sig;
  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        init_contents_busy_sig <= '1';
      else
        if init_contents_method = init_contents_method_S_0000 then
          init_contents_busy_sig <= '0';
        elsif init_contents_method = init_contents_method_S_0001 then
          init_contents_busy_sig <= tmp_0031;
        end if;
      end if;
    end if;
  end process;

  init_contents_req_sig <= init_contents_req;
  ready_contents_return <= ready_contents_return_sig;
  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        ready_contents_return_sig <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0158 then
          ready_contents_return_sig <= binary_expr_00189;
        end if;
      end if;
    end if;
  end process;

  ready_contents_busy <= ready_contents_busy_sig;
  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        ready_contents_busy_sig <= '1';
      else
        if ready_contents_method = ready_contents_method_S_0000 then
          ready_contents_busy_sig <= '0';
        elsif ready_contents_method = ready_contents_method_S_0001 then
          ready_contents_busy_sig <= tmp_0118;
        end if;
      end if;
    end if;
  end process;

  ready_contents_req_sig <= ready_contents_req;
  action_return <= action_return_sig;
  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        action_return_sig <= (others => '0');
      else
        if action_method = action_method_S_0080 then
          action_return_sig <= action_v_0204;
        end if;
      end if;
    end if;
  end process;

  action_busy <= action_busy_sig;
  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        action_busy_sig <= '1';
      else
        if action_method = action_method_S_0000 then
          action_busy_sig <= '0';
        elsif action_method = action_method_S_0001 then
          action_busy_sig <= tmp_0219;
        end if;
      end if;
    end if;
  end process;

  action_req_sig <= action_req;

  -- expressions
  tmp_0001 <= arg0_in_sig when arg0_we_sig = '1' else class_arg0_0010;
  tmp_0002 <= arg1_in_sig when arg1_we_sig = '1' else class_arg1_0011;
  tmp_0003 <= init_contents_req_local or init_contents_req_sig;
  tmp_0004 <= ready_contents_req_local or ready_contents_req_sig;
  tmp_0005 <= action_req_local or action_req_sig;
  tmp_0006 <= not pack_req_flag_d;
  tmp_0007 <= pack_req_flag and tmp_0006;
  tmp_0008 <= pack_req_flag or pack_req_flag_d;
  tmp_0009 <= pack_req_flag or pack_req_flag_d;
  tmp_0010 <= '1' when pack_method /= pack_method_S_0000 else '0';
  tmp_0011 <= '1' when pack_method /= pack_method_S_0001 else '0';
  tmp_0012 <= tmp_0011 and pack_req_flag_edge;
  tmp_0013 <= tmp_0010 and tmp_0012;
  tmp_0014 <= (32-1 downto 16 => pack_a_0012(15)) & pack_a_0012;
  tmp_0015 <= (32-1 downto 16 => pack_b_0013(15)) & pack_b_0013;
  tmp_0016 <= (32-1 downto 16 => pack_c_0014(15)) & pack_c_0014;
  tmp_0017 <= (32-1 downto 16 => pack_d_0015(15)) & pack_d_0015;
  tmp_0018 <= signed(tmp_0014) and X"000000ff";
  tmp_0019 <= signed(tmp_0015) and X"000000ff";
  tmp_0020 <= signed(tmp_0016) and X"000000ff";
  tmp_0021 <= signed(tmp_0017) and X"000000ff";
  tmp_0022 <= tmp_0018(7 downto 0) & (24-1 downto 0 => '0');
  tmp_0023 <= tmp_0019(15 downto 0) & (16-1 downto 0 => '0');
  tmp_0024 <= tmp_0020(23 downto 0) & (8-1 downto 0 => '0');
  tmp_0025 <= tmp_0022 + tmp_0023;
  tmp_0026 <= tmp_0025 + tmp_0024;
  tmp_0027 <= tmp_0026 + tmp_0021;
  tmp_0028 <= not init_contents_req_flag_d;
  tmp_0029 <= init_contents_req_flag and tmp_0028;
  tmp_0030 <= init_contents_req_flag or init_contents_req_flag_d;
  tmp_0031 <= init_contents_req_flag or init_contents_req_flag_d;
  tmp_0032 <= '1' when pack_busy = '0' else '0';
  tmp_0033 <= '1' when pack_req_local = '0' else '0';
  tmp_0034 <= tmp_0032 and tmp_0033;
  tmp_0035 <= '1' when tmp_0034 = '1' else '0';
  tmp_0036 <= '1' when pack_busy = '0' else '0';
  tmp_0037 <= '1' when pack_req_local = '0' else '0';
  tmp_0038 <= tmp_0036 and tmp_0037;
  tmp_0039 <= '1' when tmp_0038 = '1' else '0';
  tmp_0040 <= '1' when pack_busy = '0' else '0';
  tmp_0041 <= '1' when pack_req_local = '0' else '0';
  tmp_0042 <= tmp_0040 and tmp_0041;
  tmp_0043 <= '1' when tmp_0042 = '1' else '0';
  tmp_0044 <= '1' when pack_busy = '0' else '0';
  tmp_0045 <= '1' when pack_req_local = '0' else '0';
  tmp_0046 <= tmp_0044 and tmp_0045;
  tmp_0047 <= '1' when tmp_0046 = '1' else '0';
  tmp_0048 <= '1' when pack_busy = '0' else '0';
  tmp_0049 <= '1' when pack_req_local = '0' else '0';
  tmp_0050 <= tmp_0048 and tmp_0049;
  tmp_0051 <= '1' when tmp_0050 = '1' else '0';
  tmp_0052 <= '1' when pack_busy = '0' else '0';
  tmp_0053 <= '1' when pack_req_local = '0' else '0';
  tmp_0054 <= tmp_0052 and tmp_0053;
  tmp_0055 <= '1' when tmp_0054 = '1' else '0';
  tmp_0056 <= '1' when pack_busy = '0' else '0';
  tmp_0057 <= '1' when pack_req_local = '0' else '0';
  tmp_0058 <= tmp_0056 and tmp_0057;
  tmp_0059 <= '1' when tmp_0058 = '1' else '0';
  tmp_0060 <= '1' when pack_busy = '0' else '0';
  tmp_0061 <= '1' when pack_req_local = '0' else '0';
  tmp_0062 <= tmp_0060 and tmp_0061;
  tmp_0063 <= '1' when tmp_0062 = '1' else '0';
  tmp_0064 <= '1' when pack_busy = '0' else '0';
  tmp_0065 <= '1' when pack_req_local = '0' else '0';
  tmp_0066 <= tmp_0064 and tmp_0065;
  tmp_0067 <= '1' when tmp_0066 = '1' else '0';
  tmp_0068 <= '1' when pack_busy = '0' else '0';
  tmp_0069 <= '1' when pack_req_local = '0' else '0';
  tmp_0070 <= tmp_0068 and tmp_0069;
  tmp_0071 <= '1' when tmp_0070 = '1' else '0';
  tmp_0072 <= '1' when class_misc_0008_simple_div_busy = '0' else '0';
  tmp_0073 <= '1' when class_misc_0008_simple_div_req = '0' else '0';
  tmp_0074 <= tmp_0072 and tmp_0073;
  tmp_0075 <= '1' when tmp_0074 = '1' else '0';
  tmp_0076 <= '1' when class_misc_0008_simple_div_busy = '0' else '0';
  tmp_0077 <= '1' when class_misc_0008_simple_div_req = '0' else '0';
  tmp_0078 <= tmp_0076 and tmp_0077;
  tmp_0079 <= '1' when tmp_0078 = '1' else '0';
  tmp_0080 <= '1' when binary_expr_00061 = '1' else '0';
  tmp_0081 <= '1' when binary_expr_00061 = '0' else '0';
  tmp_0082 <= '1' when class_misc_0008_i_to_4digit_ascii_busy = '0' else '0';
  tmp_0083 <= '1' when class_misc_0008_i_to_4digit_ascii_req = '0' else '0';
  tmp_0084 <= tmp_0082 and tmp_0083;
  tmp_0085 <= '1' when tmp_0084 = '1' else '0';
  tmp_0086 <= '1' when class_misc_0008_i_to_4digit_ascii_busy = '0' else '0';
  tmp_0087 <= '1' when class_misc_0008_i_to_4digit_ascii_req = '0' else '0';
  tmp_0088 <= tmp_0086 and tmp_0087;
  tmp_0089 <= '1' when tmp_0088 = '1' else '0';
  tmp_0090 <= '1' when class_misc_0008_i_to_4digit_ascii_busy = '0' else '0';
  tmp_0091 <= '1' when class_misc_0008_i_to_4digit_ascii_req = '0' else '0';
  tmp_0092 <= tmp_0090 and tmp_0091;
  tmp_0093 <= '1' when tmp_0092 = '1' else '0';
  tmp_0094 <= '1' when binary_expr_00065 = '1' else '0';
  tmp_0095 <= '1' when binary_expr_00065 = '0' else '0';
  tmp_0096 <= '1' when class_misc_0008_i_to_4digit_ascii_busy = '0' else '0';
  tmp_0097 <= '1' when class_misc_0008_i_to_4digit_ascii_req = '0' else '0';
  tmp_0098 <= tmp_0096 and tmp_0097;
  tmp_0099 <= '1' when tmp_0098 = '1' else '0';
  tmp_0100 <= '1' when class_misc_0008_i_to_4digit_ascii_busy = '0' else '0';
  tmp_0101 <= '1' when class_misc_0008_i_to_4digit_ascii_req = '0' else '0';
  tmp_0102 <= tmp_0100 and tmp_0101;
  tmp_0103 <= '1' when tmp_0102 = '1' else '0';
  tmp_0104 <= '1' when class_misc_0008_i_to_4digit_ascii_busy = '0' else '0';
  tmp_0105 <= '1' when class_misc_0008_i_to_4digit_ascii_req = '0' else '0';
  tmp_0106 <= tmp_0104 and tmp_0105;
  tmp_0107 <= '1' when tmp_0106 = '1' else '0';
  tmp_0108 <= '1' when init_contents_method /= init_contents_method_S_0000 else '0';
  tmp_0109 <= '1' when init_contents_method /= init_contents_method_S_0001 else '0';
  tmp_0110 <= tmp_0109 and init_contents_req_flag_edge;
  tmp_0111 <= tmp_0108 and tmp_0110;
  tmp_0112 <= X"00000028";
  tmp_0113 <= '1' when init_contents_bytes_2_0053 > X"00000000" else '0';
  tmp_0114 <= '1' when init_contents_bytes_1_0057 > X"00000000" else '0';
  tmp_0115 <= not ready_contents_req_flag_d;
  tmp_0116 <= ready_contents_req_flag and tmp_0115;
  tmp_0117 <= ready_contents_req_flag or ready_contents_req_flag_d;
  tmp_0118 <= ready_contents_req_flag or ready_contents_req_flag_d;
  tmp_0119 <= '1' when binary_expr_00071 = '1' else '0';
  tmp_0120 <= '1' when binary_expr_00071 = '0' else '0';
  tmp_0121 <= '1' when binary_expr_00159 = '1' else '0';
  tmp_0122 <= '1' when binary_expr_00159 = '0' else '0';
  tmp_0123 <= '1' when binary_expr_00182 = '1' else '0';
  tmp_0124 <= '1' when binary_expr_00182 = '0' else '0';
  tmp_0125 <= '1' when ready_contents_method /= ready_contents_method_S_0000 else '0';
  tmp_0126 <= '1' when ready_contents_method /= ready_contents_method_S_0001 else '0';
  tmp_0127 <= tmp_0126 and ready_contents_req_flag_edge;
  tmp_0128 <= tmp_0125 and tmp_0127;
  tmp_0129 <= '1' when ready_contents_i_0069 < field_access_00070 else '0';
  tmp_0130 <= ready_contents_i_0069 + X"00000001";
  tmp_0131 <= ready_contents_i_0069(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0132 <= tmp_0131 + X"00000000";
  tmp_0133 <= (24-1 downto 0 => ready_contents_v_0073(31)) & ready_contents_v_0073(31 downto 24);
  tmp_0134 <= ready_contents_i_0069(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0135 <= tmp_0133(32 - 24 - 1 downto 0);
  tmp_0136 <= tmp_0134 + X"00000001";
  tmp_0137 <= (16-1 downto 0 => ready_contents_v_0073(31)) & ready_contents_v_0073(31 downto 16);
  tmp_0138 <= ready_contents_i_0069(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0139 <= tmp_0137(32 - 24 - 1 downto 0);
  tmp_0140 <= tmp_0138 + X"00000002";
  tmp_0141 <= (8-1 downto 0 => ready_contents_v_0073(31)) & ready_contents_v_0073(31 downto 8);
  tmp_0142 <= ready_contents_i_0069(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0143 <= tmp_0141(32 - 24 - 1 downto 0);
  tmp_0144 <= tmp_0142 + X"00000003";
  tmp_0145 <= ready_contents_v_0073;
  tmp_0146 <= tmp_0145(32 - 24 - 1 downto 0);
  tmp_0147 <= X"00000020";
  tmp_0148 <= tmp_0147 + X"00000000";
  tmp_0149 <= (24-1 downto 0 => class_content_length_field_2_0007(31)) & class_content_length_field_2_0007(31 downto 24);
  tmp_0150 <= X"00000020";
  tmp_0151 <= tmp_0149(32 - 24 - 1 downto 0);
  tmp_0152 <= tmp_0150 + X"00000001";
  tmp_0153 <= (16-1 downto 0 => class_content_length_field_2_0007(31)) & class_content_length_field_2_0007(31 downto 16);
  tmp_0154 <= X"00000020";
  tmp_0155 <= tmp_0153(32 - 24 - 1 downto 0);
  tmp_0156 <= tmp_0154 + X"00000002";
  tmp_0157 <= (8-1 downto 0 => class_content_length_field_2_0007(31)) & class_content_length_field_2_0007(31 downto 8);
  tmp_0158 <= X"00000020";
  tmp_0159 <= tmp_0157(32 - 24 - 1 downto 0);
  tmp_0160 <= tmp_0158 + X"00000003";
  tmp_0161 <= class_content_length_field_2_0007;
  tmp_0162 <= X"00000024";
  tmp_0163 <= tmp_0161(32 - 24 - 1 downto 0);
  tmp_0164 <= tmp_0162 + X"00000000";
  tmp_0165 <= (24-1 downto 0 => class_content_length_field_1_0006(31)) & class_content_length_field_1_0006(31 downto 24);
  tmp_0166 <= X"00000024";
  tmp_0167 <= tmp_0165(32 - 24 - 1 downto 0);
  tmp_0168 <= tmp_0166 + X"00000001";
  tmp_0169 <= (16-1 downto 0 => class_content_length_field_1_0006(31)) & class_content_length_field_1_0006(31 downto 16);
  tmp_0170 <= X"00000024";
  tmp_0171 <= tmp_0169(32 - 24 - 1 downto 0);
  tmp_0172 <= tmp_0170 + X"00000002";
  tmp_0173 <= (8-1 downto 0 => class_content_length_field_1_0006(31)) & class_content_length_field_1_0006(31 downto 8);
  tmp_0174 <= X"00000024";
  tmp_0175 <= tmp_0173(32 - 24 - 1 downto 0);
  tmp_0176 <= tmp_0174 + X"00000003";
  tmp_0177 <= class_content_length_field_1_0006;
  tmp_0178 <= X"00000028";
  tmp_0179 <= tmp_0177(32 - 24 - 1 downto 0);
  tmp_0180 <= tmp_0178 + X"00000000";
  tmp_0181 <= (24-1 downto 0 => class_content_length_field_0_0005(31)) & class_content_length_field_0_0005(31 downto 24);
  tmp_0182 <= X"00000028";
  tmp_0183 <= tmp_0181(32 - 24 - 1 downto 0);
  tmp_0184 <= tmp_0182 + X"00000001";
  tmp_0185 <= (16-1 downto 0 => class_content_length_field_0_0005(31)) & class_content_length_field_0_0005(31 downto 16);
  tmp_0186 <= X"00000028";
  tmp_0187 <= tmp_0185(32 - 24 - 1 downto 0);
  tmp_0188 <= tmp_0186 + X"00000002";
  tmp_0189 <= (8-1 downto 0 => class_content_length_field_0_0005(31)) & class_content_length_field_0_0005(31 downto 8);
  tmp_0190 <= X"00000028";
  tmp_0191 <= tmp_0189(32 - 24 - 1 downto 0);
  tmp_0192 <= tmp_0190 + X"00000003";
  tmp_0193 <= class_content_length_field_0_0005;
  tmp_0194 <= tmp_0193(32 - 24 - 1 downto 0);
  tmp_0195 <= '1' when ready_contents_i_0158 < class_content_words_0004 else '0';
  tmp_0196 <= ready_contents_i_0158 + X"00000001";
  tmp_0197 <= ready_contents_offset_0156 + ready_contents_i_0158;
  tmp_0198 <= tmp_0197(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0199 <= tmp_0198 + X"00000000";
  tmp_0200 <= (24-1 downto 0 => ready_contents_v_0161(31)) & ready_contents_v_0161(31 downto 24);
  tmp_0201 <= ready_contents_ptr_0163 + X"00000001";
  tmp_0202 <= tmp_0200(32 - 24 - 1 downto 0);
  tmp_0203 <= (16-1 downto 0 => ready_contents_v_0161(31)) & ready_contents_v_0161(31 downto 16);
  tmp_0204 <= ready_contents_ptr_0163 + X"00000002";
  tmp_0205 <= tmp_0203(32 - 24 - 1 downto 0);
  tmp_0206 <= (8-1 downto 0 => ready_contents_v_0161(31)) & ready_contents_v_0161(31 downto 8);
  tmp_0207 <= ready_contents_ptr_0163 + X"00000003";
  tmp_0208 <= tmp_0206(32 - 24 - 1 downto 0);
  tmp_0209 <= ready_contents_v_0161;
  tmp_0210 <= '1' when ready_contents_i_0158 = X"00000005" else '0';
  tmp_0211 <= tmp_0209(32 - 24 - 1 downto 0);
  tmp_0212 <= ready_contents_ptr_0163 + X"00000002";
  tmp_0213 <= ready_contents_ptr_0163 + X"00000003";
  tmp_0214 <= field_access_00187 + class_content_words_0004;
  tmp_0215 <= tmp_0214(29 downto 0) & (2-1 downto 0 => '0');
  tmp_0216 <= not action_req_flag_d;
  tmp_0217 <= action_req_flag and tmp_0216;
  tmp_0218 <= action_req_flag or action_req_flag_d;
  tmp_0219 <= action_req_flag or action_req_flag_d;
  tmp_0220 <= '1' when binary_expr_00195 = '1' else '0';
  tmp_0221 <= '1' when binary_expr_00195 = '0' else '0';
  tmp_0222 <= '1' when action_S_0191 = X"00000000" else '0';
  tmp_0223 <= '1' when action_S_0191 = X"00000001" else '0';
  tmp_0224 <= '1' when action_S_0191 = X"00000002" else '0';
  tmp_0225 <= '1' when action_S_0191 = X"00000003" else '0';
  tmp_0226 <= '1' when action_S_0191 = X"00000004" else '0';
  tmp_0227 <= '1' when action_S_0191 = X"00000005" else '0';
  tmp_0228 <= '1' when class_misc_0008_isHex_busy = '0' else '0';
  tmp_0229 <= '1' when class_misc_0008_isHex_req = '0' else '0';
  tmp_0230 <= tmp_0228 and tmp_0229;
  tmp_0231 <= '1' when tmp_0230 = '1' else '0';
  tmp_0232 <= '1' when method_result_00199 = '1' else '0';
  tmp_0233 <= '1' when method_result_00199 = '0' else '0';
  tmp_0234 <= '1' when class_misc_0008_isHex_busy = '0' else '0';
  tmp_0235 <= '1' when class_misc_0008_isHex_req = '0' else '0';
  tmp_0236 <= tmp_0234 and tmp_0235;
  tmp_0237 <= '1' when tmp_0236 = '1' else '0';
  tmp_0238 <= '1' when method_result_00200 = '1' else '0';
  tmp_0239 <= '1' when method_result_00200 = '0' else '0';
  tmp_0240 <= '1' when binary_expr_00201 = '1' else '0';
  tmp_0241 <= '1' when binary_expr_00201 = '0' else '0';
  tmp_0242 <= '1' when binary_expr_00202 = '1' else '0';
  tmp_0243 <= '1' when binary_expr_00202 = '0' else '0';
  tmp_0244 <= '1' when binary_expr_00203 = '1' else '0';
  tmp_0245 <= '1' when binary_expr_00203 = '0' else '0';
  tmp_0246 <= '1' when binary_expr_00205 = '1' else '0';
  tmp_0247 <= '1' when binary_expr_00205 = '0' else '0';
  tmp_0248 <= '1' when class_misc_0008_toHex2_busy = '0' else '0';
  tmp_0249 <= '1' when class_misc_0008_toHex2_req = '0' else '0';
  tmp_0250 <= tmp_0248 and tmp_0249;
  tmp_0251 <= '1' when tmp_0250 = '1' else '0';
  tmp_0252 <= '1' when action_method /= action_method_S_0000 else '0';
  tmp_0253 <= '1' when action_method /= action_method_S_0001 else '0';
  tmp_0254 <= tmp_0253 and action_req_flag_edge;
  tmp_0255 <= tmp_0252 and tmp_0254;
  tmp_0256 <= action_len_sig when action_req_sig = '1' else action_len_local;
  tmp_0257 <= '1' when action_i_0194 < action_len_0190 else '0';
  tmp_0258 <= action_i_0194 + X"00000001";
  tmp_0259 <= '1' when action_b_0197 = X"3d" else '0';
  tmp_0260 <= '1' when action_b_0197 = X"76" else '0';
  tmp_0261 <= '1' when action_b_0197 = X"3f" else '0';
  tmp_0262 <= '1' when action_S_0191 = X"00000005" else '0';

  -- sequencers
  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_method <= pack_method_IDLE;
        pack_method_delay <= (others => '0');
      else
        case (pack_method) is
          when pack_method_IDLE => 
            pack_method <= pack_method_S_0000;
          when pack_method_S_0000 => 
            pack_method <= pack_method_S_0001;
          when pack_method_S_0001 => 
            if tmp_0008 = '1' then
              pack_method <= pack_method_S_0002;
            end if;
          when pack_method_S_0002 => 
            pack_method <= pack_method_S_0016;
          when pack_method_S_0016 => 
            pack_method <= pack_method_S_0000;
          when pack_method_S_0017 => 
            pack_method <= pack_method_S_0000;
          when others => null;
        end case;
        pack_req_flag_d <= pack_req_flag;
        if (tmp_0010 and tmp_0012) = '1' then
          pack_method <= pack_method_S_0001;
        end if;
      end if;
    end if;
  end process;

  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        init_contents_method <= init_contents_method_IDLE;
        init_contents_method_delay <= (others => '0');
      else
        case (init_contents_method) is
          when init_contents_method_IDLE => 
            init_contents_method <= init_contents_method_S_0000;
          when init_contents_method_S_0000 => 
            init_contents_method <= init_contents_method_S_0001;
          when init_contents_method_S_0001 => 
            if tmp_0030 = '1' then
              init_contents_method <= init_contents_method_S_0002;
            end if;
          when init_contents_method_S_0002 => 
            init_contents_method <= init_contents_method_S_0003;
          when init_contents_method_S_0003 => 
            init_contents_method <= init_contents_method_S_0003_body;
          when init_contents_method_S_0004 => 
            init_contents_method <= init_contents_method_S_0005;
          when init_contents_method_S_0005 => 
            init_contents_method <= init_contents_method_S_0006;
          when init_contents_method_S_0006 => 
            init_contents_method <= init_contents_method_S_0006_body;
          when init_contents_method_S_0007 => 
            init_contents_method <= init_contents_method_S_0008;
          when init_contents_method_S_0008 => 
            init_contents_method <= init_contents_method_S_0009;
          when init_contents_method_S_0009 => 
            init_contents_method <= init_contents_method_S_0009_body;
          when init_contents_method_S_0010 => 
            init_contents_method <= init_contents_method_S_0011;
          when init_contents_method_S_0011 => 
            init_contents_method <= init_contents_method_S_0012;
          when init_contents_method_S_0012 => 
            init_contents_method <= init_contents_method_S_0012_body;
          when init_contents_method_S_0013 => 
            init_contents_method <= init_contents_method_S_0014;
          when init_contents_method_S_0014 => 
            init_contents_method <= init_contents_method_S_0015;
          when init_contents_method_S_0015 => 
            init_contents_method <= init_contents_method_S_0015_body;
          when init_contents_method_S_0016 => 
            init_contents_method <= init_contents_method_S_0017;
          when init_contents_method_S_0017 => 
            init_contents_method <= init_contents_method_S_0018;
          when init_contents_method_S_0018 => 
            init_contents_method <= init_contents_method_S_0018_body;
          when init_contents_method_S_0019 => 
            init_contents_method <= init_contents_method_S_0020;
          when init_contents_method_S_0020 => 
            init_contents_method <= init_contents_method_S_0021;
          when init_contents_method_S_0021 => 
            init_contents_method <= init_contents_method_S_0021_body;
          when init_contents_method_S_0022 => 
            init_contents_method <= init_contents_method_S_0023;
          when init_contents_method_S_0023 => 
            init_contents_method <= init_contents_method_S_0024;
          when init_contents_method_S_0024 => 
            init_contents_method <= init_contents_method_S_0024_body;
          when init_contents_method_S_0025 => 
            init_contents_method <= init_contents_method_S_0026;
          when init_contents_method_S_0026 => 
            init_contents_method <= init_contents_method_S_0027;
          when init_contents_method_S_0027 => 
            init_contents_method <= init_contents_method_S_0027_body;
          when init_contents_method_S_0028 => 
            init_contents_method <= init_contents_method_S_0029;
          when init_contents_method_S_0029 => 
            init_contents_method <= init_contents_method_S_0030;
          when init_contents_method_S_0030 => 
            init_contents_method <= init_contents_method_S_0030_body;
          when init_contents_method_S_0031 => 
            init_contents_method <= init_contents_method_S_0035;
          when init_contents_method_S_0035 => 
            init_contents_method <= init_contents_method_S_0035_body;
          when init_contents_method_S_0036 => 
            init_contents_method <= init_contents_method_S_0037;
          when init_contents_method_S_0037 => 
            init_contents_method <= init_contents_method_S_0038;
          when init_contents_method_S_0038 => 
            init_contents_method <= init_contents_method_S_0039;
          when init_contents_method_S_0039 => 
            init_contents_method <= init_contents_method_S_0040;
          when init_contents_method_S_0040 => 
            init_contents_method <= init_contents_method_S_0040_body;
          when init_contents_method_S_0041 => 
            init_contents_method <= init_contents_method_S_0042;
          when init_contents_method_S_0042 => 
            init_contents_method <= init_contents_method_S_0043;
          when init_contents_method_S_0043 => 
            init_contents_method <= init_contents_method_S_0044;
          when init_contents_method_S_0044 => 
            init_contents_method <= init_contents_method_S_0046;
          when init_contents_method_S_0046 => 
            if tmp_0080 = '1' then
              init_contents_method <= init_contents_method_S_0048;
            elsif tmp_0081 = '1' then
              init_contents_method <= init_contents_method_S_0055;
            end if;
          when init_contents_method_S_0047 => 
            init_contents_method <= init_contents_method_S_0070;
          when init_contents_method_S_0048 => 
            init_contents_method <= init_contents_method_S_0048_body;
          when init_contents_method_S_0049 => 
            init_contents_method <= init_contents_method_S_0050;
          when init_contents_method_S_0050 => 
            init_contents_method <= init_contents_method_S_0050_body;
          when init_contents_method_S_0051 => 
            init_contents_method <= init_contents_method_S_0052;
          when init_contents_method_S_0052 => 
            init_contents_method <= init_contents_method_S_0052_body;
          when init_contents_method_S_0053 => 
            init_contents_method <= init_contents_method_S_0054;
          when init_contents_method_S_0054 => 
            init_contents_method <= init_contents_method_S_0047;
          when init_contents_method_S_0055 => 
            init_contents_method <= init_contents_method_S_0056;
          when init_contents_method_S_0056 => 
            if tmp_0094 = '1' then
              init_contents_method <= init_contents_method_S_0058;
            elsif tmp_0095 = '1' then
              init_contents_method <= init_contents_method_S_0064;
            end if;
          when init_contents_method_S_0057 => 
            init_contents_method <= init_contents_method_S_0069;
          when init_contents_method_S_0058 => 
            init_contents_method <= init_contents_method_S_0059;
          when init_contents_method_S_0059 => 
            init_contents_method <= init_contents_method_S_0059_body;
          when init_contents_method_S_0060 => 
            init_contents_method <= init_contents_method_S_0061;
          when init_contents_method_S_0061 => 
            init_contents_method <= init_contents_method_S_0061_body;
          when init_contents_method_S_0062 => 
            init_contents_method <= init_contents_method_S_0063;
          when init_contents_method_S_0063 => 
            init_contents_method <= init_contents_method_S_0057;
          when init_contents_method_S_0064 => 
            init_contents_method <= init_contents_method_S_0066;
          when init_contents_method_S_0066 => 
            init_contents_method <= init_contents_method_S_0066_body;
          when init_contents_method_S_0067 => 
            init_contents_method <= init_contents_method_S_0068;
          when init_contents_method_S_0068 => 
            init_contents_method <= init_contents_method_S_0057;
          when init_contents_method_S_0069 => 
            init_contents_method <= init_contents_method_S_0047;
          when init_contents_method_S_0070 => 
            init_contents_method <= init_contents_method_S_0000;
          when init_contents_method_S_0003_body => 
            init_contents_method <= init_contents_method_S_0003_wait;
          when init_contents_method_S_0003_wait => 
            if pack_call_flag_0003 = '1' then
              init_contents_method <= init_contents_method_S_0004;
            end if;
          when init_contents_method_S_0006_body => 
            init_contents_method <= init_contents_method_S_0006_wait;
          when init_contents_method_S_0006_wait => 
            if pack_call_flag_0006 = '1' then
              init_contents_method <= init_contents_method_S_0007;
            end if;
          when init_contents_method_S_0009_body => 
            init_contents_method <= init_contents_method_S_0009_wait;
          when init_contents_method_S_0009_wait => 
            if pack_call_flag_0009 = '1' then
              init_contents_method <= init_contents_method_S_0010;
            end if;
          when init_contents_method_S_0012_body => 
            init_contents_method <= init_contents_method_S_0012_wait;
          when init_contents_method_S_0012_wait => 
            if pack_call_flag_0012 = '1' then
              init_contents_method <= init_contents_method_S_0013;
            end if;
          when init_contents_method_S_0015_body => 
            init_contents_method <= init_contents_method_S_0015_wait;
          when init_contents_method_S_0015_wait => 
            if pack_call_flag_0015 = '1' then
              init_contents_method <= init_contents_method_S_0016;
            end if;
          when init_contents_method_S_0018_body => 
            init_contents_method <= init_contents_method_S_0018_wait;
          when init_contents_method_S_0018_wait => 
            if pack_call_flag_0018 = '1' then
              init_contents_method <= init_contents_method_S_0019;
            end if;
          when init_contents_method_S_0021_body => 
            init_contents_method <= init_contents_method_S_0021_wait;
          when init_contents_method_S_0021_wait => 
            if pack_call_flag_0021 = '1' then
              init_contents_method <= init_contents_method_S_0022;
            end if;
          when init_contents_method_S_0024_body => 
            init_contents_method <= init_contents_method_S_0024_wait;
          when init_contents_method_S_0024_wait => 
            if pack_call_flag_0024 = '1' then
              init_contents_method <= init_contents_method_S_0025;
            end if;
          when init_contents_method_S_0027_body => 
            init_contents_method <= init_contents_method_S_0027_wait;
          when init_contents_method_S_0027_wait => 
            if pack_call_flag_0027 = '1' then
              init_contents_method <= init_contents_method_S_0028;
            end if;
          when init_contents_method_S_0030_body => 
            init_contents_method <= init_contents_method_S_0030_wait;
          when init_contents_method_S_0030_wait => 
            if pack_call_flag_0030 = '1' then
              init_contents_method <= init_contents_method_S_0031;
            end if;
          when init_contents_method_S_0035_body => 
            init_contents_method <= init_contents_method_S_0035_wait;
          when init_contents_method_S_0035_wait => 
            if simple_div_ext_call_flag_0035 = '1' then
              init_contents_method <= init_contents_method_S_0036;
            end if;
          when init_contents_method_S_0040_body => 
            init_contents_method <= init_contents_method_S_0040_wait;
          when init_contents_method_S_0040_wait => 
            if simple_div_ext_call_flag_0040 = '1' then
              init_contents_method <= init_contents_method_S_0041;
            end if;
          when init_contents_method_S_0048_body => 
            init_contents_method <= init_contents_method_S_0048_wait;
          when init_contents_method_S_0048_wait => 
            if i_to_4digit_ascii_ext_call_flag_0048 = '1' then
              init_contents_method <= init_contents_method_S_0049;
            end if;
          when init_contents_method_S_0050_body => 
            init_contents_method <= init_contents_method_S_0050_wait;
          when init_contents_method_S_0050_wait => 
            if i_to_4digit_ascii_ext_call_flag_0050 = '1' then
              init_contents_method <= init_contents_method_S_0051;
            end if;
          when init_contents_method_S_0052_body => 
            init_contents_method <= init_contents_method_S_0052_wait;
          when init_contents_method_S_0052_wait => 
            if i_to_4digit_ascii_ext_call_flag_0052 = '1' then
              init_contents_method <= init_contents_method_S_0053;
            end if;
          when init_contents_method_S_0059_body => 
            init_contents_method <= init_contents_method_S_0059_wait;
          when init_contents_method_S_0059_wait => 
            if i_to_4digit_ascii_ext_call_flag_0059 = '1' then
              init_contents_method <= init_contents_method_S_0060;
            end if;
          when init_contents_method_S_0061_body => 
            init_contents_method <= init_contents_method_S_0061_wait;
          when init_contents_method_S_0061_wait => 
            if i_to_4digit_ascii_ext_call_flag_0061 = '1' then
              init_contents_method <= init_contents_method_S_0062;
            end if;
          when init_contents_method_S_0066_body => 
            init_contents_method <= init_contents_method_S_0066_wait;
          when init_contents_method_S_0066_wait => 
            if i_to_4digit_ascii_ext_call_flag_0066 = '1' then
              init_contents_method <= init_contents_method_S_0067;
            end if;
          when others => null;
        end case;
        init_contents_req_flag_d <= init_contents_req_flag;
        if (tmp_0108 and tmp_0110) = '1' then
          init_contents_method <= init_contents_method_S_0001;
        end if;
      end if;
    end if;
  end process;

  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        ready_contents_method <= ready_contents_method_IDLE;
        ready_contents_method_delay <= (others => '0');
      else
        case (ready_contents_method) is
          when ready_contents_method_IDLE => 
            ready_contents_method <= ready_contents_method_S_0000;
          when ready_contents_method_S_0000 => 
            ready_contents_method <= ready_contents_method_S_0001;
          when ready_contents_method_S_0001 => 
            if tmp_0117 = '1' then
              ready_contents_method <= ready_contents_method_S_0002;
            end if;
          when ready_contents_method_S_0002 => 
            ready_contents_method <= ready_contents_method_S_0003;
          when ready_contents_method_S_0003 => 
            ready_contents_method <= ready_contents_method_S_0004;
          when ready_contents_method_S_0004 => 
            ready_contents_method <= ready_contents_method_S_0005;
          when ready_contents_method_S_0005 => 
            if tmp_0119 = '1' then
              ready_contents_method <= ready_contents_method_S_0010;
            elsif tmp_0120 = '1' then
              ready_contents_method <= ready_contents_method_S_0006;
            end if;
          when ready_contents_method_S_0006 => 
            ready_contents_method <= ready_contents_method_S_0038;
          when ready_contents_method_S_0007 => 
            ready_contents_method <= ready_contents_method_S_0009;
          when ready_contents_method_S_0009 => 
            ready_contents_method <= ready_contents_method_S_0003;
          when ready_contents_method_S_0010 => 
            ready_contents_method <= ready_contents_method_S_0011;
          when ready_contents_method_S_0011 => 
            if ready_contents_method_delay >= 2 then
              ready_contents_method_delay <= (others => '0');
              ready_contents_method <= ready_contents_method_S_0012;
            else
              ready_contents_method_delay <= ready_contents_method_delay + 1;
            end if;
          when ready_contents_method_S_0012 => 
            ready_contents_method <= ready_contents_method_S_0015;
          when ready_contents_method_S_0015 => 
            ready_contents_method <= ready_contents_method_S_0016;
          when ready_contents_method_S_0016 => 
            ready_contents_method <= ready_contents_method_S_0021;
          when ready_contents_method_S_0021 => 
            ready_contents_method <= ready_contents_method_S_0022;
          when ready_contents_method_S_0022 => 
            ready_contents_method <= ready_contents_method_S_0027;
          when ready_contents_method_S_0027 => 
            ready_contents_method <= ready_contents_method_S_0028;
          when ready_contents_method_S_0028 => 
            ready_contents_method <= ready_contents_method_S_0033;
          when ready_contents_method_S_0033 => 
            ready_contents_method <= ready_contents_method_S_0034;
          when ready_contents_method_S_0034 => 
            ready_contents_method <= ready_contents_method_S_0037;
          when ready_contents_method_S_0037 => 
            ready_contents_method <= ready_contents_method_S_0007;
          when ready_contents_method_S_0038 => 
            ready_contents_method <= ready_contents_method_S_0040;
          when ready_contents_method_S_0040 => 
            ready_contents_method <= ready_contents_method_S_0041;
          when ready_contents_method_S_0041 => 
            ready_contents_method <= ready_contents_method_S_0046;
          when ready_contents_method_S_0046 => 
            ready_contents_method <= ready_contents_method_S_0047;
          when ready_contents_method_S_0047 => 
            ready_contents_method <= ready_contents_method_S_0052;
          when ready_contents_method_S_0052 => 
            ready_contents_method <= ready_contents_method_S_0053;
          when ready_contents_method_S_0053 => 
            ready_contents_method <= ready_contents_method_S_0058;
          when ready_contents_method_S_0058 => 
            ready_contents_method <= ready_contents_method_S_0059;
          when ready_contents_method_S_0059 => 
            ready_contents_method <= ready_contents_method_S_0064;
          when ready_contents_method_S_0064 => 
            ready_contents_method <= ready_contents_method_S_0065;
          when ready_contents_method_S_0065 => 
            ready_contents_method <= ready_contents_method_S_0070;
          when ready_contents_method_S_0070 => 
            ready_contents_method <= ready_contents_method_S_0071;
          when ready_contents_method_S_0071 => 
            ready_contents_method <= ready_contents_method_S_0076;
          when ready_contents_method_S_0076 => 
            ready_contents_method <= ready_contents_method_S_0077;
          when ready_contents_method_S_0077 => 
            ready_contents_method <= ready_contents_method_S_0082;
          when ready_contents_method_S_0082 => 
            ready_contents_method <= ready_contents_method_S_0083;
          when ready_contents_method_S_0083 => 
            ready_contents_method <= ready_contents_method_S_0088;
          when ready_contents_method_S_0088 => 
            ready_contents_method <= ready_contents_method_S_0089;
          when ready_contents_method_S_0089 => 
            ready_contents_method <= ready_contents_method_S_0094;
          when ready_contents_method_S_0094 => 
            ready_contents_method <= ready_contents_method_S_0095;
          when ready_contents_method_S_0095 => 
            ready_contents_method <= ready_contents_method_S_0100;
          when ready_contents_method_S_0100 => 
            ready_contents_method <= ready_contents_method_S_0101;
          when ready_contents_method_S_0101 => 
            ready_contents_method <= ready_contents_method_S_0106;
          when ready_contents_method_S_0106 => 
            ready_contents_method <= ready_contents_method_S_0107;
          when ready_contents_method_S_0107 => 
            ready_contents_method <= ready_contents_method_S_0110;
          when ready_contents_method_S_0110 => 
            ready_contents_method <= ready_contents_method_S_0111;
          when ready_contents_method_S_0111 => 
            ready_contents_method <= ready_contents_method_S_0113;
          when ready_contents_method_S_0113 => 
            ready_contents_method <= ready_contents_method_S_0114;
          when ready_contents_method_S_0114 => 
            if tmp_0121 = '1' then
              ready_contents_method <= ready_contents_method_S_0119;
            elsif tmp_0122 = '1' then
              ready_contents_method <= ready_contents_method_S_0115;
            end if;
          when ready_contents_method_S_0115 => 
            ready_contents_method <= ready_contents_method_S_0155;
          when ready_contents_method_S_0116 => 
            ready_contents_method <= ready_contents_method_S_0118;
          when ready_contents_method_S_0118 => 
            ready_contents_method <= ready_contents_method_S_0113;
          when ready_contents_method_S_0119 => 
            if ready_contents_method_delay >= 2 then
              ready_contents_method_delay <= (others => '0');
              ready_contents_method <= ready_contents_method_S_0120;
            else
              ready_contents_method_delay <= ready_contents_method_delay + 1;
            end if;
          when ready_contents_method_S_0120 => 
            ready_contents_method <= ready_contents_method_S_0125;
          when ready_contents_method_S_0125 => 
            ready_contents_method <= ready_contents_method_S_0126;
          when ready_contents_method_S_0126 => 
            ready_contents_method <= ready_contents_method_S_0130;
          when ready_contents_method_S_0130 => 
            ready_contents_method <= ready_contents_method_S_0131;
          when ready_contents_method_S_0131 => 
            ready_contents_method <= ready_contents_method_S_0135;
          when ready_contents_method_S_0135 => 
            ready_contents_method <= ready_contents_method_S_0136;
          when ready_contents_method_S_0136 => 
            ready_contents_method <= ready_contents_method_S_0140;
          when ready_contents_method_S_0140 => 
            ready_contents_method <= ready_contents_method_S_0141;
          when ready_contents_method_S_0141 => 
            ready_contents_method <= ready_contents_method_S_0145;
          when ready_contents_method_S_0145 => 
            if tmp_0123 = '1' then
              ready_contents_method <= ready_contents_method_S_0147;
            elsif tmp_0124 = '1' then
              ready_contents_method <= ready_contents_method_S_0146;
            end if;
          when ready_contents_method_S_0146 => 
            ready_contents_method <= ready_contents_method_S_0154;
          when ready_contents_method_S_0147 => 
            ready_contents_method <= ready_contents_method_S_0148;
          when ready_contents_method_S_0148 => 
            ready_contents_method <= ready_contents_method_S_0150;
          when ready_contents_method_S_0150 => 
            ready_contents_method <= ready_contents_method_S_0151;
          when ready_contents_method_S_0151 => 
            ready_contents_method <= ready_contents_method_S_0153;
          when ready_contents_method_S_0153 => 
            ready_contents_method <= ready_contents_method_S_0146;
          when ready_contents_method_S_0154 => 
            ready_contents_method <= ready_contents_method_S_0116;
          when ready_contents_method_S_0155 => 
            ready_contents_method <= ready_contents_method_S_0156;
          when ready_contents_method_S_0156 => 
            ready_contents_method <= ready_contents_method_S_0158;
          when ready_contents_method_S_0158 => 
            ready_contents_method <= ready_contents_method_S_0000;
          when ready_contents_method_S_0159 => 
            ready_contents_method <= ready_contents_method_S_0000;
          when others => null;
        end case;
        ready_contents_req_flag_d <= ready_contents_req_flag;
        if (tmp_0125 and tmp_0127) = '1' then
          ready_contents_method <= ready_contents_method_S_0001;
        end if;
      end if;
    end if;
  end process;

  process (clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        action_method <= action_method_IDLE;
        action_method_delay <= (others => '0');
      else
        case (action_method) is
          when action_method_IDLE => 
            action_method <= action_method_S_0000;
          when action_method_S_0000 => 
            action_method <= action_method_S_0001;
          when action_method_S_0001 => 
            if tmp_0218 = '1' then
              action_method <= action_method_S_0002;
            end if;
          when action_method_S_0002 => 
            action_method <= action_method_S_0006;
          when action_method_S_0006 => 
            action_method <= action_method_S_0007;
          when action_method_S_0007 => 
            if tmp_0220 = '1' then
              action_method <= action_method_S_0012;
            elsif tmp_0221 = '1' then
              action_method <= action_method_S_0008;
            end if;
          when action_method_S_0008 => 
            action_method <= action_method_S_0068;
          when action_method_S_0009 => 
            action_method <= action_method_S_0011;
          when action_method_S_0011 => 
            action_method <= action_method_S_0006;
          when action_method_S_0012 => 
            if action_method_delay >= 2 then
              action_method_delay <= (others => '0');
              action_method <= action_method_S_0013;
            else
              action_method_delay <= action_method_delay + 1;
            end if;
          when action_method_S_0013 => 
            action_method <= action_method_S_0014;
          when action_method_S_0014 => 
            if tmp_0222 = '1' then
              action_method <= action_method_S_0058;
            elsif tmp_0223 = '1' then
              action_method <= action_method_S_0049;
            elsif tmp_0224 = '1' then
              action_method <= action_method_S_0040;
            elsif tmp_0225 = '1' then
              action_method <= action_method_S_0030;
            elsif tmp_0226 = '1' then
              action_method <= action_method_S_0020;
            elsif tmp_0227 = '1' then
              action_method <= action_method_S_0018;
            else
              action_method <= action_method_S_0016;
            end if;
          when action_method_S_0015 => 
            action_method <= action_method_S_0067;
          when action_method_S_0016 => 
            action_method <= action_method_S_0017;
          when action_method_S_0017 => 
            action_method <= action_method_S_0015;
          when action_method_S_0018 => 
            action_method <= action_method_S_0015;
          when action_method_S_0019 => 
            action_method <= action_method_S_0016;
          when action_method_S_0020 => 
            action_method <= action_method_S_0020_body;
          when action_method_S_0021 => 
            if tmp_0232 = '1' then
              action_method <= action_method_S_0023;
            elsif tmp_0233 = '1' then
              action_method <= action_method_S_0026;
            end if;
          when action_method_S_0022 => 
            action_method <= action_method_S_0028;
          when action_method_S_0023 => 
            action_method <= action_method_S_0025;
          when action_method_S_0025 => 
            action_method <= action_method_S_0022;
          when action_method_S_0026 => 
            action_method <= action_method_S_0027;
          when action_method_S_0027 => 
            action_method <= action_method_S_0022;
          when action_method_S_0028 => 
            action_method <= action_method_S_0015;
          when action_method_S_0029 => 
            action_method <= action_method_S_0018;
          when action_method_S_0030 => 
            action_method <= action_method_S_0030_body;
          when action_method_S_0031 => 
            if tmp_0238 = '1' then
              action_method <= action_method_S_0033;
            elsif tmp_0239 = '1' then
              action_method <= action_method_S_0036;
            end if;
          when action_method_S_0032 => 
            action_method <= action_method_S_0038;
          when action_method_S_0033 => 
            action_method <= action_method_S_0035;
          when action_method_S_0035 => 
            action_method <= action_method_S_0032;
          when action_method_S_0036 => 
            action_method <= action_method_S_0037;
          when action_method_S_0037 => 
            action_method <= action_method_S_0032;
          when action_method_S_0038 => 
            action_method <= action_method_S_0015;
          when action_method_S_0039 => 
            action_method <= action_method_S_0020;
          when action_method_S_0040 => 
            action_method <= action_method_S_0041;
          when action_method_S_0041 => 
            if tmp_0240 = '1' then
              action_method <= action_method_S_0043;
            elsif tmp_0241 = '1' then
              action_method <= action_method_S_0045;
            end if;
          when action_method_S_0042 => 
            action_method <= action_method_S_0047;
          when action_method_S_0043 => 
            action_method <= action_method_S_0044;
          when action_method_S_0044 => 
            action_method <= action_method_S_0042;
          when action_method_S_0045 => 
            action_method <= action_method_S_0046;
          when action_method_S_0046 => 
            action_method <= action_method_S_0042;
          when action_method_S_0047 => 
            action_method <= action_method_S_0015;
          when action_method_S_0048 => 
            action_method <= action_method_S_0030;
          when action_method_S_0049 => 
            action_method <= action_method_S_0050;
          when action_method_S_0050 => 
            if tmp_0242 = '1' then
              action_method <= action_method_S_0052;
            elsif tmp_0243 = '1' then
              action_method <= action_method_S_0054;
            end if;
          when action_method_S_0051 => 
            action_method <= action_method_S_0056;
          when action_method_S_0052 => 
            action_method <= action_method_S_0053;
          when action_method_S_0053 => 
            action_method <= action_method_S_0051;
          when action_method_S_0054 => 
            action_method <= action_method_S_0055;
          when action_method_S_0055 => 
            action_method <= action_method_S_0051;
          when action_method_S_0056 => 
            action_method <= action_method_S_0015;
          when action_method_S_0057 => 
            action_method <= action_method_S_0040;
          when action_method_S_0058 => 
            action_method <= action_method_S_0059;
          when action_method_S_0059 => 
            if tmp_0244 = '1' then
              action_method <= action_method_S_0061;
            elsif tmp_0245 = '1' then
              action_method <= action_method_S_0063;
            end if;
          when action_method_S_0060 => 
            action_method <= action_method_S_0065;
          when action_method_S_0061 => 
            action_method <= action_method_S_0062;
          when action_method_S_0062 => 
            action_method <= action_method_S_0060;
          when action_method_S_0063 => 
            action_method <= action_method_S_0064;
          when action_method_S_0064 => 
            action_method <= action_method_S_0060;
          when action_method_S_0065 => 
            action_method <= action_method_S_0015;
          when action_method_S_0066 => 
            action_method <= action_method_S_0049;
          when action_method_S_0067 => 
            action_method <= action_method_S_0009;
          when action_method_S_0068 => 
            action_method <= action_method_S_0070;
          when action_method_S_0070 => 
            if tmp_0246 = '1' then
              action_method <= action_method_S_0072;
            elsif tmp_0247 = '1' then
              action_method <= action_method_S_0077;
            end if;
          when action_method_S_0071 => 
            action_method <= action_method_S_0080;
          when action_method_S_0072 => 
            action_method <= action_method_S_0072_body;
          when action_method_S_0073 => 
            action_method <= action_method_S_0076;
          when action_method_S_0076 => 
            action_method <= action_method_S_0071;
          when action_method_S_0077 => 
            action_method <= action_method_S_0079;
          when action_method_S_0079 => 
            action_method <= action_method_S_0071;
          when action_method_S_0080 => 
            action_method <= action_method_S_0000;
          when action_method_S_0081 => 
            action_method <= action_method_S_0000;
          when action_method_S_0020_body => 
            action_method <= action_method_S_0020_wait;
          when action_method_S_0020_wait => 
            if isHex_ext_call_flag_0020 = '1' then
              action_method <= action_method_S_0021;
            end if;
          when action_method_S_0030_body => 
            action_method <= action_method_S_0030_wait;
          when action_method_S_0030_wait => 
            if isHex_ext_call_flag_0030 = '1' then
              action_method <= action_method_S_0031;
            end if;
          when action_method_S_0072_body => 
            action_method <= action_method_S_0072_wait;
          when action_method_S_0072_wait => 
            if toHex2_ext_call_flag_0072 = '1' then
              action_method <= action_method_S_0073;
            end if;
          when others => null;
        end case;
        action_req_flag_d <= action_req_flag;
        if (tmp_0252 and tmp_0254) = '1' then
          action_method <= action_method_S_0001;
        end if;
      end if;
    end if;
  end process;


  class_resp_0000_clk <= clk_sig;

  class_resp_0000_reset <= reset_sig;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_resp_0000_data_address <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0011 and ready_contents_method_delay = 0 then
          class_resp_0000_data_address <= ready_contents_i_0069;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_resp_0000_data_oe <= '0';
      else
        if ready_contents_method = ready_contents_method_S_0011 and ready_contents_method_delay = 0 then
          class_resp_0000_data_oe <= '1';
        else
          class_resp_0000_data_oe <= '0';
        end if;
      end if;
    end if;
  end process;

  class_buffer_0002_clk <= clk_sig;

  class_buffer_0002_reset <= reset_sig;

  class_buffer_0002_address <= buffer_address_sig;

  class_buffer_0002_din <= buffer_din_sig;

  class_buffer_0002_we <= buffer_we_sig;

  class_buffer_0002_oe <= buffer_oe_sig;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_buffer_0002_address_b <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0015 then
          class_buffer_0002_address_b <= binary_expr_00077;
        elsif ready_contents_method = ready_contents_method_S_0021 then
          class_buffer_0002_address_b <= binary_expr_00082;
        elsif ready_contents_method = ready_contents_method_S_0027 then
          class_buffer_0002_address_b <= binary_expr_00087;
        elsif ready_contents_method = ready_contents_method_S_0033 then
          class_buffer_0002_address_b <= binary_expr_00092;
        elsif ready_contents_method = ready_contents_method_S_0040 then
          class_buffer_0002_address_b <= binary_expr_00097;
        elsif ready_contents_method = ready_contents_method_S_0046 then
          class_buffer_0002_address_b <= binary_expr_00102;
        elsif ready_contents_method = ready_contents_method_S_0052 then
          class_buffer_0002_address_b <= binary_expr_00107;
        elsif ready_contents_method = ready_contents_method_S_0058 then
          class_buffer_0002_address_b <= binary_expr_00112;
        elsif ready_contents_method = ready_contents_method_S_0064 then
          class_buffer_0002_address_b <= binary_expr_00117;
        elsif ready_contents_method = ready_contents_method_S_0070 then
          class_buffer_0002_address_b <= binary_expr_00122;
        elsif ready_contents_method = ready_contents_method_S_0076 then
          class_buffer_0002_address_b <= binary_expr_00127;
        elsif ready_contents_method = ready_contents_method_S_0082 then
          class_buffer_0002_address_b <= binary_expr_00132;
        elsif ready_contents_method = ready_contents_method_S_0088 then
          class_buffer_0002_address_b <= binary_expr_00137;
        elsif ready_contents_method = ready_contents_method_S_0094 then
          class_buffer_0002_address_b <= binary_expr_00142;
        elsif ready_contents_method = ready_contents_method_S_0100 then
          class_buffer_0002_address_b <= binary_expr_00147;
        elsif ready_contents_method = ready_contents_method_S_0106 then
          class_buffer_0002_address_b <= binary_expr_00152;
        elsif ready_contents_method = ready_contents_method_S_0125 then
          class_buffer_0002_address_b <= binary_expr_00166;
        elsif ready_contents_method = ready_contents_method_S_0130 then
          class_buffer_0002_address_b <= binary_expr_00170;
        elsif ready_contents_method = ready_contents_method_S_0135 then
          class_buffer_0002_address_b <= binary_expr_00174;
        elsif ready_contents_method = ready_contents_method_S_0140 then
          class_buffer_0002_address_b <= binary_expr_00178;
        elsif ready_contents_method = ready_contents_method_S_0148 then
          class_buffer_0002_address_b <= binary_expr_00183;
        elsif ready_contents_method = ready_contents_method_S_0151 then
          class_buffer_0002_address_b <= binary_expr_00185;
        elsif action_method = action_method_S_0012 and action_method_delay = 0 then
          class_buffer_0002_address_b <= action_i_0194;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_buffer_0002_din_b <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0016 then
          class_buffer_0002_din_b <= tmp_0135;
        elsif ready_contents_method = ready_contents_method_S_0022 then
          class_buffer_0002_din_b <= tmp_0139;
        elsif ready_contents_method = ready_contents_method_S_0028 then
          class_buffer_0002_din_b <= tmp_0143;
        elsif ready_contents_method = ready_contents_method_S_0034 then
          class_buffer_0002_din_b <= tmp_0146;
        elsif ready_contents_method = ready_contents_method_S_0041 then
          class_buffer_0002_din_b <= tmp_0151;
        elsif ready_contents_method = ready_contents_method_S_0047 then
          class_buffer_0002_din_b <= tmp_0155;
        elsif ready_contents_method = ready_contents_method_S_0053 then
          class_buffer_0002_din_b <= tmp_0159;
        elsif ready_contents_method = ready_contents_method_S_0059 then
          class_buffer_0002_din_b <= tmp_0163;
        elsif ready_contents_method = ready_contents_method_S_0065 then
          class_buffer_0002_din_b <= tmp_0167;
        elsif ready_contents_method = ready_contents_method_S_0071 then
          class_buffer_0002_din_b <= tmp_0171;
        elsif ready_contents_method = ready_contents_method_S_0077 then
          class_buffer_0002_din_b <= tmp_0175;
        elsif ready_contents_method = ready_contents_method_S_0083 then
          class_buffer_0002_din_b <= tmp_0179;
        elsif ready_contents_method = ready_contents_method_S_0089 then
          class_buffer_0002_din_b <= tmp_0183;
        elsif ready_contents_method = ready_contents_method_S_0095 then
          class_buffer_0002_din_b <= tmp_0187;
        elsif ready_contents_method = ready_contents_method_S_0101 then
          class_buffer_0002_din_b <= tmp_0191;
        elsif ready_contents_method = ready_contents_method_S_0107 then
          class_buffer_0002_din_b <= tmp_0194;
        elsif ready_contents_method = ready_contents_method_S_0126 then
          class_buffer_0002_din_b <= tmp_0202;
        elsif ready_contents_method = ready_contents_method_S_0131 then
          class_buffer_0002_din_b <= tmp_0205;
        elsif ready_contents_method = ready_contents_method_S_0136 then
          class_buffer_0002_din_b <= tmp_0208;
        elsif ready_contents_method = ready_contents_method_S_0141 then
          class_buffer_0002_din_b <= tmp_0211;
        elsif ready_contents_method = ready_contents_method_S_0148 then
          class_buffer_0002_din_b <= class_arg0_0010;
        elsif ready_contents_method = ready_contents_method_S_0151 then
          class_buffer_0002_din_b <= class_arg1_0011;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_buffer_0002_we_b <= '0';
      else
        if ready_contents_method = ready_contents_method_S_0016 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0022 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0028 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0034 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0041 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0047 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0053 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0059 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0065 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0071 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0077 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0083 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0089 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0095 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0101 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0107 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0126 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0131 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0136 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0141 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0148 then
          class_buffer_0002_we_b <= '1';
        elsif ready_contents_method = ready_contents_method_S_0151 then
          class_buffer_0002_we_b <= '1';
        else
          class_buffer_0002_we_b <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_buffer_0002_oe_b <= '0';
      else
        if action_method = action_method_S_0012 and action_method_delay = 0 then
          class_buffer_0002_oe_b <= '1';
        else
          class_buffer_0002_oe_b <= '0';
        end if;
      end if;
    end if;
  end process;

  class_data_0003_clk <= clk_sig;

  class_data_0003_reset <= reset_sig;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_data_0003_address_b <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0002 then
          class_data_0003_address_b <= X"00000000";
        elsif init_contents_method = init_contents_method_S_0005 then
          class_data_0003_address_b <= X"00000001";
        elsif init_contents_method = init_contents_method_S_0008 then
          class_data_0003_address_b <= X"00000002";
        elsif init_contents_method = init_contents_method_S_0011 then
          class_data_0003_address_b <= X"00000003";
        elsif init_contents_method = init_contents_method_S_0014 then
          class_data_0003_address_b <= X"00000004";
        elsif init_contents_method = init_contents_method_S_0017 then
          class_data_0003_address_b <= X"00000005";
        elsif init_contents_method = init_contents_method_S_0020 then
          class_data_0003_address_b <= X"00000006";
        elsif init_contents_method = init_contents_method_S_0023 then
          class_data_0003_address_b <= X"00000007";
        elsif init_contents_method = init_contents_method_S_0026 then
          class_data_0003_address_b <= X"00000008";
        elsif init_contents_method = init_contents_method_S_0029 then
          class_data_0003_address_b <= X"00000009";
        elsif ready_contents_method = ready_contents_method_S_0119 and ready_contents_method_delay = 0 then
          class_data_0003_address_b <= ready_contents_i_0158;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_data_0003_din_b <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0004 then
          class_data_0003_din_b <= method_result_00031;
        elsif init_contents_method = init_contents_method_S_0007 then
          class_data_0003_din_b <= method_result_00033;
        elsif init_contents_method = init_contents_method_S_0010 then
          class_data_0003_din_b <= method_result_00035;
        elsif init_contents_method = init_contents_method_S_0013 then
          class_data_0003_din_b <= method_result_00037;
        elsif init_contents_method = init_contents_method_S_0016 then
          class_data_0003_din_b <= method_result_00039;
        elsif init_contents_method = init_contents_method_S_0019 then
          class_data_0003_din_b <= method_result_00041;
        elsif init_contents_method = init_contents_method_S_0022 then
          class_data_0003_din_b <= method_result_00043;
        elsif init_contents_method = init_contents_method_S_0025 then
          class_data_0003_din_b <= method_result_00045;
        elsif init_contents_method = init_contents_method_S_0028 then
          class_data_0003_din_b <= method_result_00047;
        elsif init_contents_method = init_contents_method_S_0031 then
          class_data_0003_din_b <= method_result_00049;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_data_0003_we_b <= '0';
      else
        if init_contents_method = init_contents_method_S_0004 then
          class_data_0003_we_b <= '1';
        elsif init_contents_method = init_contents_method_S_0007 then
          class_data_0003_we_b <= '1';
        elsif init_contents_method = init_contents_method_S_0010 then
          class_data_0003_we_b <= '1';
        elsif init_contents_method = init_contents_method_S_0013 then
          class_data_0003_we_b <= '1';
        elsif init_contents_method = init_contents_method_S_0016 then
          class_data_0003_we_b <= '1';
        elsif init_contents_method = init_contents_method_S_0019 then
          class_data_0003_we_b <= '1';
        elsif init_contents_method = init_contents_method_S_0022 then
          class_data_0003_we_b <= '1';
        elsif init_contents_method = init_contents_method_S_0025 then
          class_data_0003_we_b <= '1';
        elsif init_contents_method = init_contents_method_S_0028 then
          class_data_0003_we_b <= '1';
        elsif init_contents_method = init_contents_method_S_0031 then
          class_data_0003_we_b <= '1';
        else
          class_data_0003_we_b <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_data_0003_oe_b <= '0';
      else
        if ready_contents_method = ready_contents_method_S_0119 and ready_contents_method_delay = 0 then
          class_data_0003_oe_b <= '1';
        else
          class_data_0003_oe_b <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_content_words_0004 <= X"00000008";
      else
        if init_contents_method = init_contents_method_S_0031 then
          class_content_words_0004 <= X"0000000a";
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_content_length_field_0_0005 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0053 then
          class_content_length_field_0_0005 <= method_result_00064;
        elsif init_contents_method = init_contents_method_S_0062 then
          class_content_length_field_0_0005 <= method_result_00067;
        elsif init_contents_method = init_contents_method_S_0067 then
          class_content_length_field_0_0005 <= method_result_00068;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_content_length_field_1_0006 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0051 then
          class_content_length_field_1_0006 <= method_result_00063;
        elsif init_contents_method = init_contents_method_S_0060 then
          class_content_length_field_1_0006 <= method_result_00066;
        elsif init_contents_method = init_contents_method_S_0064 then
          class_content_length_field_1_0006 <= X"20202020";
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_content_length_field_2_0007 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0049 then
          class_content_length_field_2_0007 <= method_result_00062;
        elsif init_contents_method = init_contents_method_S_0058 then
          class_content_length_field_2_0007 <= X"20202020";
        elsif init_contents_method = init_contents_method_S_0064 then
          class_content_length_field_2_0007 <= X"20202020";
        end if;
      end if;
    end if;
  end process;

  class_misc_0008_clk <= clk_sig;

  class_misc_0008_reset <= reset_sig;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_simple_div_n <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0035_body and init_contents_method_delay = 0 then
          class_misc_0008_simple_div_n <= init_contents_v_0050;
        elsif init_contents_method = init_contents_method_S_0040_body and init_contents_method_delay = 0 then
          class_misc_0008_simple_div_n <= init_contents_v_0050;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_simple_div_d <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0035_body and init_contents_method_delay = 0 then
          class_misc_0008_simple_div_d <= X"05f5e100";
        elsif init_contents_method = init_contents_method_S_0040_body and init_contents_method_delay = 0 then
          class_misc_0008_simple_div_d <= X"00002710";
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_i_to_4digit_ascii_x <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0048_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_x <= init_contents_bytes_2_0053;
        elsif init_contents_method = init_contents_method_S_0050_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_x <= init_contents_bytes_1_0057;
        elsif init_contents_method = init_contents_method_S_0052_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_x <= init_contents_bytes_0_0059;
        elsif init_contents_method = init_contents_method_S_0059_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_x <= init_contents_bytes_1_0057;
        elsif init_contents_method = init_contents_method_S_0061_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_x <= init_contents_bytes_0_0059;
        elsif init_contents_method = init_contents_method_S_0066_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_x <= init_contents_bytes_0_0059;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_i_to_4digit_ascii_flag <= '0';
      else
        if init_contents_method = init_contents_method_S_0048_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_flag <= '0';
        elsif init_contents_method = init_contents_method_S_0050_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_flag <= '1';
        elsif init_contents_method = init_contents_method_S_0052_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_flag <= '1';
        elsif init_contents_method = init_contents_method_S_0059_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_flag <= '0';
        elsif init_contents_method = init_contents_method_S_0061_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_flag <= '1';
        elsif init_contents_method = init_contents_method_S_0066_body and init_contents_method_delay = 0 then
          class_misc_0008_i_to_4digit_ascii_flag <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_isHex_v <= (others => '0');
      else
        if action_method = action_method_S_0020_body and action_method_delay = 0 then
          class_misc_0008_isHex_v <= action_b_0197;
        elsif action_method = action_method_S_0030_body and action_method_delay = 0 then
          class_misc_0008_isHex_v <= action_b_0197;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_toHex2_v0 <= (others => '0');
      else
        if action_method = action_method_S_0072_body and action_method_delay = 0 then
          class_misc_0008_toHex2_v0 <= action_v0_0192;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_toHex2_v1 <= (others => '0');
      else
        if action_method = action_method_S_0072_body and action_method_delay = 0 then
          class_misc_0008_toHex2_v1 <= action_v1_0193;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_simple_div_req <= '0';
      else
        if init_contents_method = init_contents_method_S_0035_body then
          class_misc_0008_simple_div_req <= '1';
        elsif init_contents_method = init_contents_method_S_0040_body then
          class_misc_0008_simple_div_req <= '1';
        else
          class_misc_0008_simple_div_req <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_i_to_4digit_ascii_req <= '0';
      else
        if init_contents_method = init_contents_method_S_0048_body then
          class_misc_0008_i_to_4digit_ascii_req <= '1';
        elsif init_contents_method = init_contents_method_S_0050_body then
          class_misc_0008_i_to_4digit_ascii_req <= '1';
        elsif init_contents_method = init_contents_method_S_0052_body then
          class_misc_0008_i_to_4digit_ascii_req <= '1';
        elsif init_contents_method = init_contents_method_S_0059_body then
          class_misc_0008_i_to_4digit_ascii_req <= '1';
        elsif init_contents_method = init_contents_method_S_0061_body then
          class_misc_0008_i_to_4digit_ascii_req <= '1';
        elsif init_contents_method = init_contents_method_S_0066_body then
          class_misc_0008_i_to_4digit_ascii_req <= '1';
        else
          class_misc_0008_i_to_4digit_ascii_req <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_isHex_req <= '0';
      else
        if action_method = action_method_S_0020_body then
          class_misc_0008_isHex_req <= '1';
        elsif action_method = action_method_S_0030_body then
          class_misc_0008_isHex_req <= '1';
        else
          class_misc_0008_isHex_req <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_misc_0008_toHex2_req <= '0';
      else
        if action_method = action_method_S_0072_body then
          class_misc_0008_toHex2_req <= '1';
        else
          class_misc_0008_toHex2_req <= '0';
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_arg0_0010 <= X"20";
      else
        if action_method = action_method_S_0073 then
          class_arg0_0010 <= action_v0_0192;
        elsif action_method = action_method_S_0077 then
          class_arg0_0010 <= X"3f";
        else
          class_arg0_0010 <= class_arg0_0010_mux;
        end if;
      end if;
    end if;
  end process;

  class_arg0_0010_mux <= tmp_0001;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        class_arg1_0011 <= X"20";
      else
        if action_method = action_method_S_0073 then
          class_arg1_0011 <= action_v1_0193;
        elsif action_method = action_method_S_0077 then
          class_arg1_0011 <= X"3f";
        else
          class_arg1_0011 <= class_arg1_0011_mux;
        end if;
      end if;
    end if;
  end process;

  class_arg1_0011_mux <= tmp_0002;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_a_0012 <= (others => '0');
      else
        if pack_method = pack_method_S_0001 then
          pack_a_0012 <= pack_a_local;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_a_local <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0003_body and init_contents_method_delay = 0 then
          pack_a_local <= X"003c";
        elsif init_contents_method = init_contents_method_S_0006_body and init_contents_method_delay = 0 then
          pack_a_local <= X"006c";
        elsif init_contents_method = init_contents_method_S_0009_body and init_contents_method_delay = 0 then
          pack_a_local <= X"006f";
        elsif init_contents_method = init_contents_method_S_0012_body and init_contents_method_delay = 0 then
          pack_a_local <= X"0041";
        elsif init_contents_method = init_contents_method_S_0015_body and init_contents_method_delay = 0 then
          pack_a_local <= X"006d";
        elsif init_contents_method = init_contents_method_S_0018_body and init_contents_method_delay = 0 then
          pack_a_local <= X"003f";
        elsif init_contents_method = init_contents_method_S_0021_body and init_contents_method_delay = 0 then
          pack_a_local <= X"003c";
        elsif init_contents_method = init_contents_method_S_0024_body and init_contents_method_delay = 0 then
          pack_a_local <= X"0064";
        elsif init_contents_method = init_contents_method_S_0027_body and init_contents_method_delay = 0 then
          pack_a_local <= X"002f";
        elsif init_contents_method = init_contents_method_S_0030_body and init_contents_method_delay = 0 then
          pack_a_local <= X"006c";
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_b_0013 <= (others => '0');
      else
        if pack_method = pack_method_S_0001 then
          pack_b_0013 <= pack_b_local;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_b_local <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0003_body and init_contents_method_delay = 0 then
          pack_b_local <= X"0068";
        elsif init_contents_method = init_contents_method_S_0006_body and init_contents_method_delay = 0 then
          pack_b_local <= X"003e";
        elsif init_contents_method = init_contents_method_S_0009_body and init_contents_method_delay = 0 then
          pack_b_local <= X"0064";
        elsif init_contents_method = init_contents_method_S_0012_body and init_contents_method_delay = 0 then
          pack_b_local <= X"0072";
        elsif init_contents_method = init_contents_method_S_0015_body and init_contents_method_delay = 0 then
          pack_b_local <= X"0065";
        elsif init_contents_method = init_contents_method_S_0018_body and init_contents_method_delay = 0 then
          pack_b_local <= X"003d";
        elsif init_contents_method = init_contents_method_S_0021_body and init_contents_method_delay = 0 then
          pack_b_local <= X"002f";
        elsif init_contents_method = init_contents_method_S_0024_body and init_contents_method_delay = 0 then
          pack_b_local <= X"0079";
        elsif init_contents_method = init_contents_method_S_0027_body and init_contents_method_delay = 0 then
          pack_b_local <= X"0068";
        elsif init_contents_method = init_contents_method_S_0030_body and init_contents_method_delay = 0 then
          pack_b_local <= X"003e";
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_c_0014 <= (others => '0');
      else
        if pack_method = pack_method_S_0001 then
          pack_c_0014 <= pack_c_local;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_c_local <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0003_body and init_contents_method_delay = 0 then
          pack_c_local <= X"0074";
        elsif init_contents_method = init_contents_method_S_0006_body and init_contents_method_delay = 0 then
          pack_c_local <= X"003c";
        elsif init_contents_method = init_contents_method_S_0009_body and init_contents_method_delay = 0 then
          pack_c_local <= X"0079";
        elsif init_contents_method = init_contents_method_S_0012_body and init_contents_method_delay = 0 then
          pack_c_local <= X"0067";
        elsif init_contents_method = init_contents_method_S_0015_body and init_contents_method_delay = 0 then
          pack_c_local <= X"006e";
        elsif init_contents_method = init_contents_method_S_0018_body and init_contents_method_delay = 0 then
          pack_c_local <= X"0020";
        elsif init_contents_method = init_contents_method_S_0021_body and init_contents_method_delay = 0 then
          pack_c_local <= X"0062";
        elsif init_contents_method = init_contents_method_S_0024_body and init_contents_method_delay = 0 then
          pack_c_local <= X"003e";
        elsif init_contents_method = init_contents_method_S_0027_body and init_contents_method_delay = 0 then
          pack_c_local <= X"0074";
        elsif init_contents_method = init_contents_method_S_0030_body and init_contents_method_delay = 0 then
          pack_c_local <= X"000a";
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_d_0015 <= (others => '0');
      else
        if pack_method = pack_method_S_0001 then
          pack_d_0015 <= pack_d_local;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_d_local <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0003_body and init_contents_method_delay = 0 then
          pack_d_local <= X"006d";
        elsif init_contents_method = init_contents_method_S_0006_body and init_contents_method_delay = 0 then
          pack_d_local <= X"0062";
        elsif init_contents_method = init_contents_method_S_0009_body and init_contents_method_delay = 0 then
          pack_d_local <= X"003e";
        elsif init_contents_method = init_contents_method_S_0012_body and init_contents_method_delay = 0 then
          pack_d_local <= X"0075";
        elsif init_contents_method = init_contents_method_S_0015_body and init_contents_method_delay = 0 then
          pack_d_local <= X"0074";
        elsif init_contents_method = init_contents_method_S_0018_body and init_contents_method_delay = 0 then
          pack_d_local <= X"0020";
        elsif init_contents_method = init_contents_method_S_0021_body and init_contents_method_delay = 0 then
          pack_d_local <= X"006f";
        elsif init_contents_method = init_contents_method_S_0024_body and init_contents_method_delay = 0 then
          pack_d_local <= X"003c";
        elsif init_contents_method = init_contents_method_S_0027_body and init_contents_method_delay = 0 then
          pack_d_local <= X"006d";
        elsif init_contents_method = init_contents_method_S_0030_body and init_contents_method_delay = 0 then
          pack_d_local <= X"000a";
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00016 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          cast_expr_00016 <= signed(tmp_0014);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00017 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          binary_expr_00017 <= tmp_0018;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00018 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          binary_expr_00018 <= tmp_0022;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00019 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          cast_expr_00019 <= signed(tmp_0015);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00020 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          binary_expr_00020 <= tmp_0019;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00021 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          binary_expr_00021 <= tmp_0023;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00022 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          binary_expr_00022 <= tmp_0025;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00023 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          cast_expr_00023 <= signed(tmp_0016);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00024 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          binary_expr_00024 <= tmp_0020;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00025 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          binary_expr_00025 <= tmp_0024;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00026 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          binary_expr_00026 <= tmp_0026;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00027 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          cast_expr_00027 <= signed(tmp_0017);
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00028 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          binary_expr_00028 <= tmp_0021;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00029 <= (others => '0');
      else
        if pack_method = pack_method_S_0002 then
          binary_expr_00029 <= tmp_0027;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00031 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0003_wait then
          method_result_00031 <= pack_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00033 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0006_wait then
          method_result_00033 <= pack_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00035 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0009_wait then
          method_result_00035 <= pack_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00037 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0012_wait then
          method_result_00037 <= pack_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00039 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0015_wait then
          method_result_00039 <= pack_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00041 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0018_wait then
          method_result_00041 <= pack_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00043 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0021_wait then
          method_result_00043 <= pack_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00045 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0024_wait then
          method_result_00045 <= pack_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00047 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0027_wait then
          method_result_00047 <= pack_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00049 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0030_wait then
          method_result_00049 <= pack_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        init_contents_v_0050 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0031 then
          init_contents_v_0050 <= tmp_0112;
        elsif init_contents_method = init_contents_method_S_0039 then
          init_contents_v_0050 <= field_access_00055;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00051 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0031 then
          binary_expr_00051 <= tmp_0112;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00052 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0035_wait then
          method_result_00052 <= class_misc_0008_simple_div_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        init_contents_bytes_2_0053 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0037 then
          init_contents_bytes_2_0053 <= field_access_00054;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00054 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0036 then
          field_access_00054 <= class_misc_0008_quant_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00055 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0038 then
          field_access_00055 <= class_misc_0008_remainder_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00056 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0040_wait then
          method_result_00056 <= class_misc_0008_simple_div_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        init_contents_bytes_1_0057 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0042 then
          init_contents_bytes_1_0057 <= field_access_00058;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00058 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0041 then
          field_access_00058 <= class_misc_0008_quant_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        init_contents_bytes_0_0059 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0044 then
          init_contents_bytes_0_0059 <= field_access_00060;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00060 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0043 then
          field_access_00060 <= class_misc_0008_remainder_out;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00061 <= '0';
      else
        if init_contents_method = init_contents_method_S_0044 then
          binary_expr_00061 <= tmp_0113;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00062 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0048_wait then
          method_result_00062 <= class_misc_0008_i_to_4digit_ascii_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00063 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0050_wait then
          method_result_00063 <= class_misc_0008_i_to_4digit_ascii_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00064 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0052_wait then
          method_result_00064 <= class_misc_0008_i_to_4digit_ascii_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00065 <= '0';
      else
        if init_contents_method = init_contents_method_S_0055 then
          binary_expr_00065 <= tmp_0114;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00066 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0059_wait then
          method_result_00066 <= class_misc_0008_i_to_4digit_ascii_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00067 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0061_wait then
          method_result_00067 <= class_misc_0008_i_to_4digit_ascii_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00068 <= (others => '0');
      else
        if init_contents_method = init_contents_method_S_0066_wait then
          method_result_00068 <= class_misc_0008_i_to_4digit_ascii_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00096 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0038 then
          binary_expr_00096 <= tmp_0147;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00097 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0038 then
          binary_expr_00097 <= tmp_0148;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00099 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0041 then
          binary_expr_00099 <= tmp_0149;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00100 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0041 then
          cast_expr_00100 <= tmp_0151;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00101 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0041 then
          binary_expr_00101 <= tmp_0150;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00102 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0041 then
          binary_expr_00102 <= tmp_0152;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00104 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0047 then
          binary_expr_00104 <= tmp_0153;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00105 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0047 then
          cast_expr_00105 <= tmp_0155;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00106 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0047 then
          binary_expr_00106 <= tmp_0154;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00107 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0047 then
          binary_expr_00107 <= tmp_0156;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00109 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0053 then
          binary_expr_00109 <= tmp_0157;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00110 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0053 then
          cast_expr_00110 <= tmp_0159;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00111 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0053 then
          binary_expr_00111 <= tmp_0158;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00112 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0053 then
          binary_expr_00112 <= tmp_0160;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00114 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0059 then
          binary_expr_00114 <= tmp_0161;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00115 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0059 then
          cast_expr_00115 <= tmp_0163;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00116 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0059 then
          binary_expr_00116 <= tmp_0162;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00117 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0059 then
          binary_expr_00117 <= tmp_0164;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00119 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0065 then
          binary_expr_00119 <= tmp_0165;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00120 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0065 then
          cast_expr_00120 <= tmp_0167;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00121 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0065 then
          binary_expr_00121 <= tmp_0166;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00122 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0065 then
          binary_expr_00122 <= tmp_0168;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00124 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0071 then
          binary_expr_00124 <= tmp_0169;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00125 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0071 then
          cast_expr_00125 <= tmp_0171;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00126 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0071 then
          binary_expr_00126 <= tmp_0170;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00127 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0071 then
          binary_expr_00127 <= tmp_0172;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00129 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0077 then
          binary_expr_00129 <= tmp_0173;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00130 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0077 then
          cast_expr_00130 <= tmp_0175;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00131 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0077 then
          binary_expr_00131 <= tmp_0174;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00132 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0077 then
          binary_expr_00132 <= tmp_0176;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00134 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0083 then
          binary_expr_00134 <= tmp_0177;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00135 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0083 then
          cast_expr_00135 <= tmp_0179;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00136 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0083 then
          binary_expr_00136 <= tmp_0178;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00137 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0083 then
          binary_expr_00137 <= tmp_0180;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00139 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0089 then
          binary_expr_00139 <= tmp_0181;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00140 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0089 then
          cast_expr_00140 <= tmp_0183;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00141 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0089 then
          binary_expr_00141 <= tmp_0182;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00142 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0089 then
          binary_expr_00142 <= tmp_0184;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00144 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0095 then
          binary_expr_00144 <= tmp_0185;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00145 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0095 then
          cast_expr_00145 <= tmp_0187;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00146 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0095 then
          binary_expr_00146 <= tmp_0186;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00147 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0095 then
          binary_expr_00147 <= tmp_0188;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00149 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0101 then
          binary_expr_00149 <= tmp_0189;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00150 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0101 then
          cast_expr_00150 <= tmp_0191;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00151 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0101 then
          binary_expr_00151 <= tmp_0190;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00152 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0101 then
          binary_expr_00152 <= tmp_0192;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00154 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0107 then
          binary_expr_00154 <= tmp_0193;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00155 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0107 then
          cast_expr_00155 <= tmp_0194;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        ready_contents_offset_0156 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0111 then
          ready_contents_offset_0156 <= field_access_00157;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00157 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0110 then
          field_access_00157 <= class_resp_0000_length;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00187 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0155 then
          field_access_00187 <= class_resp_0000_length;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00188 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0156 then
          binary_expr_00188 <= tmp_0214;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00189 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0156 then
          binary_expr_00189 <= tmp_0215;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        ready_contents_i_0069 <= X"00000000";
      else
        if ready_contents_method = ready_contents_method_S_0002 then
          ready_contents_i_0069 <= X"00000000";
        elsif ready_contents_method = ready_contents_method_S_0007 then
          ready_contents_i_0069 <= tmp_0130;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        field_access_00070 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0003 then
          field_access_00070 <= class_resp_0000_length;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00071 <= '0';
      else
        if ready_contents_method = ready_contents_method_S_0004 then
          binary_expr_00071 <= tmp_0129;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        unary_expr_00072 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0007 then
          unary_expr_00072 <= tmp_0130;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        ready_contents_v_0073 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0012 then
          ready_contents_v_0073 <= array_access_00075;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00075 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0011 and ready_contents_method_delay = 2 then
          array_access_00075 <= class_resp_0000_data_dout;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00076 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0012 then
          binary_expr_00076 <= tmp_0131;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00077 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0012 then
          binary_expr_00077 <= tmp_0132;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00079 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0016 then
          binary_expr_00079 <= tmp_0133;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00080 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0016 then
          cast_expr_00080 <= tmp_0135;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00081 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0016 then
          binary_expr_00081 <= tmp_0134;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00082 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0016 then
          binary_expr_00082 <= tmp_0136;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00084 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0022 then
          binary_expr_00084 <= tmp_0137;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00085 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0022 then
          cast_expr_00085 <= tmp_0139;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00086 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0022 then
          binary_expr_00086 <= tmp_0138;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00087 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0022 then
          binary_expr_00087 <= tmp_0140;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00089 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0028 then
          binary_expr_00089 <= tmp_0141;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00090 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0028 then
          cast_expr_00090 <= tmp_0143;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00091 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0028 then
          binary_expr_00091 <= tmp_0142;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00092 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0028 then
          binary_expr_00092 <= tmp_0144;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00094 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0034 then
          binary_expr_00094 <= tmp_0145;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00095 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0034 then
          cast_expr_00095 <= tmp_0146;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        ready_contents_i_0158 <= X"00000000";
      else
        if ready_contents_method = ready_contents_method_S_0111 then
          ready_contents_i_0158 <= X"00000000";
        elsif ready_contents_method = ready_contents_method_S_0116 then
          ready_contents_i_0158 <= tmp_0196;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00159 <= '0';
      else
        if ready_contents_method = ready_contents_method_S_0113 then
          binary_expr_00159 <= tmp_0195;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        unary_expr_00160 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0116 then
          unary_expr_00160 <= tmp_0196;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        ready_contents_v_0161 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0120 then
          ready_contents_v_0161 <= array_access_00162;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00162 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0119 and ready_contents_method_delay = 2 then
          array_access_00162 <= class_data_0003_dout_b;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        ready_contents_ptr_0163 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0120 then
          ready_contents_ptr_0163 <= tmp_0198;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00164 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0120 then
          binary_expr_00164 <= tmp_0197;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00165 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0120 then
          binary_expr_00165 <= tmp_0198;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00166 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0120 then
          binary_expr_00166 <= tmp_0199;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00168 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0126 then
          binary_expr_00168 <= tmp_0200;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00169 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0126 then
          cast_expr_00169 <= tmp_0202;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00170 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0126 then
          binary_expr_00170 <= tmp_0201;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00172 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0131 then
          binary_expr_00172 <= tmp_0203;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00173 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0131 then
          cast_expr_00173 <= tmp_0205;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00174 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0131 then
          binary_expr_00174 <= tmp_0204;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00176 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0136 then
          binary_expr_00176 <= tmp_0206;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00177 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0136 then
          cast_expr_00177 <= tmp_0208;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00178 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0136 then
          binary_expr_00178 <= tmp_0207;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00180 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0141 then
          binary_expr_00180 <= tmp_0209;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        cast_expr_00181 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0141 then
          cast_expr_00181 <= tmp_0211;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00182 <= '0';
      else
        if ready_contents_method = ready_contents_method_S_0141 then
          binary_expr_00182 <= tmp_0210;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00183 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0147 then
          binary_expr_00183 <= tmp_0212;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00185 <= (others => '0');
      else
        if ready_contents_method = ready_contents_method_S_0150 then
          binary_expr_00185 <= tmp_0213;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        action_len_0190 <= (others => '0');
      else
        if action_method = action_method_S_0001 then
          action_len_0190 <= tmp_0256;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        action_S_0191 <= X"00000000";
      else
        if action_method = action_method_S_0002 then
          action_S_0191 <= X"00000000";
        elsif action_method = action_method_S_0016 then
          action_S_0191 <= X"00000000";
        elsif action_method = action_method_S_0023 then
          action_S_0191 <= X"00000005";
        elsif action_method = action_method_S_0026 then
          action_S_0191 <= X"00000000";
        elsif action_method = action_method_S_0033 then
          action_S_0191 <= X"00000004";
        elsif action_method = action_method_S_0036 then
          action_S_0191 <= X"00000000";
        elsif action_method = action_method_S_0043 then
          action_S_0191 <= X"00000003";
        elsif action_method = action_method_S_0045 then
          action_S_0191 <= X"00000000";
        elsif action_method = action_method_S_0052 then
          action_S_0191 <= X"00000002";
        elsif action_method = action_method_S_0054 then
          action_S_0191 <= X"00000000";
        elsif action_method = action_method_S_0061 then
          action_S_0191 <= X"00000001";
        elsif action_method = action_method_S_0063 then
          action_S_0191 <= X"00000000";
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        action_v0_0192 <= X"00";
      else
        if action_method = action_method_S_0002 then
          action_v0_0192 <= X"00";
        elsif action_method = action_method_S_0033 then
          action_v0_0192 <= action_b_0197;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        action_v1_0193 <= X"00";
      else
        if action_method = action_method_S_0002 then
          action_v1_0193 <= X"00";
        elsif action_method = action_method_S_0023 then
          action_v1_0193 <= action_b_0197;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        action_v_0204 <= X"00000000";
      else
        if action_method = action_method_S_0068 then
          action_v_0204 <= X"00000000";
        elsif action_method = action_method_S_0073 then
          action_v_0204 <= method_result_00206;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00205 <= '0';
      else
        if action_method = action_method_S_0068 then
          binary_expr_00205 <= tmp_0262;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        action_i_0194 <= X"00000000";
      else
        if action_method = action_method_S_0002 then
          action_i_0194 <= X"00000000";
        elsif action_method = action_method_S_0009 then
          action_i_0194 <= tmp_0258;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00195 <= '0';
      else
        if action_method = action_method_S_0006 then
          binary_expr_00195 <= tmp_0257;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        unary_expr_00196 <= (others => '0');
      else
        if action_method = action_method_S_0009 then
          unary_expr_00196 <= tmp_0258;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        action_b_0197 <= (others => '0');
      else
        if action_method = action_method_S_0013 then
          action_b_0197 <= array_access_00198;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        array_access_00198 <= (others => '0');
      else
        if action_method = action_method_S_0012 and action_method_delay = 2 then
          array_access_00198 <= class_buffer_0002_dout_b;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00199 <= '0';
      else
        if action_method = action_method_S_0020_wait then
          method_result_00199 <= class_misc_0008_isHex_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00200 <= '0';
      else
        if action_method = action_method_S_0030_wait then
          method_result_00200 <= class_misc_0008_isHex_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00201 <= '0';
      else
        if action_method = action_method_S_0040 then
          binary_expr_00201 <= tmp_0259;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00202 <= '0';
      else
        if action_method = action_method_S_0049 then
          binary_expr_00202 <= tmp_0260;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        binary_expr_00203 <= '0';
      else
        if action_method = action_method_S_0058 then
          binary_expr_00203 <= tmp_0261;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        method_result_00206 <= (others => '0');
      else
        if action_method = action_method_S_0072_wait then
          method_result_00206 <= class_misc_0008_toHex2_return;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_return <= (others => '0');
      else
        if pack_method = pack_method_S_0016 then
          pack_return <= binary_expr_00029;
        end if;
      end if;
    end if;
  end process;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_busy <= '0';
      else
        if pack_method = pack_method_S_0000 then
          pack_busy <= '0';
        elsif pack_method = pack_method_S_0001 then
          pack_busy <= tmp_0009;
        end if;
      end if;
    end if;
  end process;

  pack_req_flag <= pack_req_local;

  process(clk)
  begin
    if clk'event and clk = '1' then
      if reset = '1' then
        pack_req_local <= '0';
      else
        if init_contents_method = init_contents_method_S_0003_body then
          pack_req_local <= '1';
        elsif init_contents_method = init_contents_method_S_0006_body then
          pack_req_local <= '1';
        elsif init_contents_method = init_contents_method_S_0009_body then
          pack_req_local <= '1';
        elsif init_contents_method = init_contents_method_S_0012_body then
          pack_req_local <= '1';
        elsif init_contents_method = init_contents_method_S_0015_body then
          pack_req_local <= '1';
        elsif init_contents_method = init_contents_method_S_0018_body then
          pack_req_local <= '1';
        elsif init_contents_method = init_contents_method_S_0021_body then
          pack_req_local <= '1';
        elsif init_contents_method = init_contents_method_S_0024_body then
          pack_req_local <= '1';
        elsif init_contents_method = init_contents_method_S_0027_body then
          pack_req_local <= '1';
        elsif init_contents_method = init_contents_method_S_0030_body then
          pack_req_local <= '1';
        else
          pack_req_local <= '0';
        end if;
      end if;
    end if;
  end process;

  init_contents_req_flag <= tmp_0003;

  ready_contents_req_flag <= tmp_0004;

  action_req_flag <= tmp_0005;

  pack_req_flag_edge <= tmp_0007;

  init_contents_req_flag_edge <= tmp_0029;

  pack_call_flag_0003 <= tmp_0035;

  pack_call_flag_0006 <= tmp_0039;

  pack_call_flag_0009 <= tmp_0043;

  pack_call_flag_0012 <= tmp_0047;

  pack_call_flag_0015 <= tmp_0051;

  pack_call_flag_0018 <= tmp_0055;

  pack_call_flag_0021 <= tmp_0059;

  pack_call_flag_0024 <= tmp_0063;

  pack_call_flag_0027 <= tmp_0067;

  pack_call_flag_0030 <= tmp_0071;

  simple_div_ext_call_flag_0035 <= tmp_0075;

  simple_div_ext_call_flag_0040 <= tmp_0079;

  i_to_4digit_ascii_ext_call_flag_0048 <= tmp_0085;

  i_to_4digit_ascii_ext_call_flag_0050 <= tmp_0089;

  i_to_4digit_ascii_ext_call_flag_0052 <= tmp_0093;

  i_to_4digit_ascii_ext_call_flag_0059 <= tmp_0099;

  i_to_4digit_ascii_ext_call_flag_0061 <= tmp_0103;

  i_to_4digit_ascii_ext_call_flag_0066 <= tmp_0107;

  ready_contents_req_flag_edge <= tmp_0116;

  action_req_flag_edge <= tmp_0217;

  isHex_ext_call_flag_0020 <= tmp_0231;

  isHex_ext_call_flag_0030 <= tmp_0237;

  toHex2_ext_call_flag_0072 <= tmp_0251;


  inst_class_resp_0000 : http_response_header
  port map(
    clk => class_resp_0000_clk,
    reset => class_resp_0000_reset,
    data_length => class_resp_0000_data_length,
    data_address => class_resp_0000_data_address,
    data_din => class_resp_0000_data_din,
    data_dout => class_resp_0000_data_dout,
    data_we => class_resp_0000_data_we,
    data_oe => class_resp_0000_data_oe,
    length => class_resp_0000_length
  );

  inst_class_buffer_0002 : dualportram
  generic map(
    WIDTH => 8,
    DEPTH => 13,
    WORDS => 8192
  )
  port map(
    clk => class_buffer_0002_clk,
    reset => class_buffer_0002_reset,
    length => class_buffer_0002_length,
    address => class_buffer_0002_address,
    din => class_buffer_0002_din,
    dout => class_buffer_0002_dout,
    we => class_buffer_0002_we,
    oe => class_buffer_0002_oe,
    address_b => class_buffer_0002_address_b,
    din_b => class_buffer_0002_din_b,
    dout_b => class_buffer_0002_dout_b,
    we_b => class_buffer_0002_we_b,
    oe_b => class_buffer_0002_oe_b
  );

  inst_class_data_0003 : singleportram
  generic map(
    WIDTH => 32,
    DEPTH => 10,
    WORDS => 1024
  )
  port map(
    clk => class_data_0003_clk,
    reset => class_data_0003_reset,
    length => class_data_0003_length,
    address_b => class_data_0003_address_b,
    din_b => class_data_0003_din_b,
    dout_b => class_data_0003_dout_b,
    we_b => class_data_0003_we_b,
    oe_b => class_data_0003_oe_b
  );

  inst_class_misc_0008 : Misc
  port map(
    clk => class_misc_0008_clk,
    reset => class_misc_0008_reset,
    quant_in => class_misc_0008_quant_in,
    quant_we => class_misc_0008_quant_we,
    quant_out => class_misc_0008_quant_out,
    remainder_in => class_misc_0008_remainder_in,
    remainder_we => class_misc_0008_remainder_we,
    remainder_out => class_misc_0008_remainder_out,
    simple_div_n => class_misc_0008_simple_div_n,
    simple_div_d => class_misc_0008_simple_div_d,
    i_to_4digit_ascii_x => class_misc_0008_i_to_4digit_ascii_x,
    i_to_4digit_ascii_flag => class_misc_0008_i_to_4digit_ascii_flag,
    isHex_v => class_misc_0008_isHex_v,
    toHex1_v => class_misc_0008_toHex1_v,
    toHex2_v0 => class_misc_0008_toHex2_v0,
    toHex2_v1 => class_misc_0008_toHex2_v1,
    simple_div_return => class_misc_0008_simple_div_return,
    simple_div_busy => class_misc_0008_simple_div_busy,
    simple_div_req => class_misc_0008_simple_div_req,
    i_to_4digit_ascii_return => class_misc_0008_i_to_4digit_ascii_return,
    i_to_4digit_ascii_busy => class_misc_0008_i_to_4digit_ascii_busy,
    i_to_4digit_ascii_req => class_misc_0008_i_to_4digit_ascii_req,
    isHex_return => class_misc_0008_isHex_return,
    isHex_busy => class_misc_0008_isHex_busy,
    isHex_req => class_misc_0008_isHex_req,
    toHex1_return => class_misc_0008_toHex1_return,
    toHex1_busy => class_misc_0008_toHex1_busy,
    toHex1_req => class_misc_0008_toHex1_req,
    toHex2_return => class_misc_0008_toHex2_return,
    toHex2_busy => class_misc_0008_toHex2_busy,
    toHex2_req => class_misc_0008_toHex2_req
  );


end RTL;
